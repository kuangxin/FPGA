//------------------------------------------------------------------------------
//   ____  ____
//  /   /\/   /
// /___/  \  /    Vendor: Xilinx
// \   \   \/     Version : 2.7
//  \   \         Application : 7 Series FPGAs Transceivers Wizard 
//  /   /         Filename : serdes_coe_init.v
// /___/   /\      
// \   \  /  \ 
//  \___\/\___\
//
//  Description : This module instantiates the modules required for
//                reset and initialisation of the Transceiver
//
// Module serdes_coe_init
// Generated by Xilinx 7 Series FPGAs Transceivers Wizard
// 
// 
// (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
// 
// This file contains confidential and proprietary information
// of Xilinx, Inc. and is protected under U.S. and
// international copyright and other intellectual property
// laws.
// 
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// Xilinx, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) Xilinx shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or Xilinx had been advised of the
// possibility of the same.
// 
// CRITICAL APPLICATIONS
// Xilinx products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of Xilinx products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
// 
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES. 


`timescale 1ns / 1ps
`define DLY #1

//***********************************Entity Declaration************************

module serdes_coe_init #
(
    parameter EXAMPLE_SIM_GTRESET_SPEEDUP            = "TRUE",                  // Simulation setting for GT SecureIP model
    parameter EXAMPLE_SIMULATION                     =  0,                      // Set to 1 for simulation
    parameter STABLE_CLOCK_PERIOD                    =  10, // Period of the stable clock driving this 
                                                                                // state-machine, unit is [ns]

    parameter EXAMPLE_USE_CHIPSCOPE                  =  0                       // Set to 1 to use Chipscope to drive resets

)
(
    input           SYSCLK_IN,
    input           SOFT_RESET_IN,
    input           DONT_RESET_ON_DATA_ERROR_IN,
    output          GT0_TX_FSM_RESET_DONE_OUT,
    output          GT0_RX_FSM_RESET_DONE_OUT,
    input           GT0_DATA_VALID_IN,
    output          GT1_TX_FSM_RESET_DONE_OUT,
    output          GT1_RX_FSM_RESET_DONE_OUT,
    input           GT1_DATA_VALID_IN,
    output          GT2_TX_FSM_RESET_DONE_OUT,
    output          GT2_RX_FSM_RESET_DONE_OUT,
    input           GT2_DATA_VALID_IN,
    output          GT3_TX_FSM_RESET_DONE_OUT,
    output          GT3_RX_FSM_RESET_DONE_OUT,
    input           GT3_DATA_VALID_IN,
    output          GT4_TX_FSM_RESET_DONE_OUT,
    output          GT4_RX_FSM_RESET_DONE_OUT,
    input           GT4_DATA_VALID_IN,
    output          GT5_TX_FSM_RESET_DONE_OUT,
    output          GT5_RX_FSM_RESET_DONE_OUT,
    input           GT5_DATA_VALID_IN,
    output          GT6_TX_FSM_RESET_DONE_OUT,
    output          GT6_RX_FSM_RESET_DONE_OUT,
    input           GT6_DATA_VALID_IN,
    output          GT7_TX_FSM_RESET_DONE_OUT,
    output          GT7_RX_FSM_RESET_DONE_OUT,
    input           GT7_DATA_VALID_IN,

    //_________________________________________________________________________
    //GT0  (X1Y0)
    //____________________________CHANNEL PORTS________________________________
    //------------------------------- CPLL Ports -------------------------------
    output          GT0_CPLLFBCLKLOST_OUT,
    output          GT0_CPLLLOCK_OUT,
    input           GT0_CPLLLOCKDETCLK_IN,
    input           GT0_CPLLRESET_IN,
    //------------------------ Channel - Clocking Ports ------------------------
    input           GT0_GTREFCLK0_IN,
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   GT0_DRPADDR_IN,
    input           GT0_DRPCLK_IN,
    input   [15:0]  GT0_DRPDI_IN,
    output  [15:0]  GT0_DRPDO_OUT,
    input           GT0_DRPEN_IN,
    output          GT0_DRPRDY_OUT,
    input           GT0_DRPWE_IN,
    //----------------------------- Loopback Ports -----------------------------
    input   [2:0]   GT0_LOOPBACK_IN,
    //------------------- RX Initialization and Reset Ports --------------------
    input           GT0_RXUSERRDY_IN,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          GT0_EYESCANDATAERROR_OUT,
    //----------------------- Receive Ports - CDR Ports ------------------------
    output          GT0_RXCDRLOCK_OUT,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           GT0_RXUSRCLK_IN,
    input           GT0_RXUSRCLK2_IN,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [15:0]  GT0_RXDATA_OUT,
    //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
    output  [1:0]   GT0_RXDISPERR_OUT,
    output  [1:0]   GT0_RXNOTINTABLE_OUT,
    //------------------------- Receive Ports - RX AFE -------------------------
    input           GT0_GTXRXP_IN,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           GT0_GTXRXN_IN,
    //---------------- Receive Ports - RX Channel Bonding Ports ----------------
    output          GT0_RXCHANBONDSEQ_OUT,
    input           GT0_RXCHBONDEN_IN,
    input   [2:0]   GT0_RXCHBONDLEVEL_IN,
    input           GT0_RXCHBONDMASTER_IN,
    output  [4:0]   GT0_RXCHBONDO_OUT,
    input           GT0_RXCHBONDSLAVE_IN,
    //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
    output          GT0_RXCHANISALIGNED_OUT,
    output          GT0_RXCHANREALIGN_OUT,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           GT0_GTRXRESET_IN,
    input           GT0_RXPMARESET_IN,
    //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    output  [1:0]   GT0_RXCHARISK_OUT,
    //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
    input   [4:0]   GT0_RXCHBONDI_IN,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          GT0_RXRESETDONE_OUT,
    //------------------- TX Initialization and Reset Ports --------------------
    input           GT0_GTTXRESET_IN,
    input           GT0_TXUSERRDY_IN,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           GT0_TXUSRCLK_IN,
    input           GT0_TXUSRCLK2_IN,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [15:0]  GT0_TXDATA_IN,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          GT0_GTXTXN_OUT,
    output          GT0_GTXTXP_OUT,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          GT0_TXOUTCLK_OUT,
    output          GT0_TXOUTCLKFABRIC_OUT,
    output          GT0_TXOUTCLKPCS_OUT,
    //------------------- Transmit Ports - TX Gearbox Ports --------------------
    input   [1:0]   GT0_TXCHARISK_IN,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    output          GT0_TXRESETDONE_OUT,

    //GT1  (X1Y1)
    //____________________________CHANNEL PORTS________________________________
    //------------------------------- CPLL Ports -------------------------------
    output          GT1_CPLLFBCLKLOST_OUT,
    output          GT1_CPLLLOCK_OUT,
    input           GT1_CPLLLOCKDETCLK_IN,
    input           GT1_CPLLRESET_IN,
    //------------------------ Channel - Clocking Ports ------------------------
    input           GT1_GTREFCLK0_IN,
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   GT1_DRPADDR_IN,
    input           GT1_DRPCLK_IN,
    input   [15:0]  GT1_DRPDI_IN,
    output  [15:0]  GT1_DRPDO_OUT,
    input           GT1_DRPEN_IN,
    output          GT1_DRPRDY_OUT,
    input           GT1_DRPWE_IN,
    //----------------------------- Loopback Ports -----------------------------
    input   [2:0]   GT1_LOOPBACK_IN,
    //------------------- RX Initialization and Reset Ports --------------------
    input           GT1_RXUSERRDY_IN,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          GT1_EYESCANDATAERROR_OUT,
    //----------------------- Receive Ports - CDR Ports ------------------------
    output          GT1_RXCDRLOCK_OUT,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           GT1_RXUSRCLK_IN,
    input           GT1_RXUSRCLK2_IN,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [15:0]  GT1_RXDATA_OUT,
    //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
    output  [1:0]   GT1_RXDISPERR_OUT,
    output  [1:0]   GT1_RXNOTINTABLE_OUT,
    //------------------------- Receive Ports - RX AFE -------------------------
    input           GT1_GTXRXP_IN,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           GT1_GTXRXN_IN,
    //---------------- Receive Ports - RX Channel Bonding Ports ----------------
    output          GT1_RXCHANBONDSEQ_OUT,
    input           GT1_RXCHBONDEN_IN,
    input   [2:0]   GT1_RXCHBONDLEVEL_IN,
    input           GT1_RXCHBONDMASTER_IN,
    output  [4:0]   GT1_RXCHBONDO_OUT,
    input           GT1_RXCHBONDSLAVE_IN,
    //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
    output          GT1_RXCHANISALIGNED_OUT,
    output          GT1_RXCHANREALIGN_OUT,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           GT1_GTRXRESET_IN,
    input           GT1_RXPMARESET_IN,
    //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    output  [1:0]   GT1_RXCHARISK_OUT,
    //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
    input   [4:0]   GT1_RXCHBONDI_IN,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          GT1_RXRESETDONE_OUT,
    //------------------- TX Initialization and Reset Ports --------------------
    input           GT1_GTTXRESET_IN,
    input           GT1_TXUSERRDY_IN,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           GT1_TXUSRCLK_IN,
    input           GT1_TXUSRCLK2_IN,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [15:0]  GT1_TXDATA_IN,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          GT1_GTXTXN_OUT,
    output          GT1_GTXTXP_OUT,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          GT1_TXOUTCLK_OUT,
    output          GT1_TXOUTCLKFABRIC_OUT,
    output          GT1_TXOUTCLKPCS_OUT,
    //------------------- Transmit Ports - TX Gearbox Ports --------------------
    input   [1:0]   GT1_TXCHARISK_IN,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    output          GT1_TXRESETDONE_OUT,

    //GT2  (X1Y2)
    //____________________________CHANNEL PORTS________________________________
    //------------------------------- CPLL Ports -------------------------------
    output          GT2_CPLLFBCLKLOST_OUT,
    output          GT2_CPLLLOCK_OUT,
    input           GT2_CPLLLOCKDETCLK_IN,
    input           GT2_CPLLRESET_IN,
    //------------------------ Channel - Clocking Ports ------------------------
    input           GT2_GTREFCLK0_IN,
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   GT2_DRPADDR_IN,
    input           GT2_DRPCLK_IN,
    input   [15:0]  GT2_DRPDI_IN,
    output  [15:0]  GT2_DRPDO_OUT,
    input           GT2_DRPEN_IN,
    output          GT2_DRPRDY_OUT,
    input           GT2_DRPWE_IN,
    //----------------------------- Loopback Ports -----------------------------
    input   [2:0]   GT2_LOOPBACK_IN,
    //------------------- RX Initialization and Reset Ports --------------------
    input           GT2_RXUSERRDY_IN,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          GT2_EYESCANDATAERROR_OUT,
    //----------------------- Receive Ports - CDR Ports ------------------------
    output          GT2_RXCDRLOCK_OUT,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           GT2_RXUSRCLK_IN,
    input           GT2_RXUSRCLK2_IN,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [15:0]  GT2_RXDATA_OUT,
    //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
    output  [1:0]   GT2_RXDISPERR_OUT,
    output  [1:0]   GT2_RXNOTINTABLE_OUT,
    //------------------------- Receive Ports - RX AFE -------------------------
    input           GT2_GTXRXP_IN,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           GT2_GTXRXN_IN,
    //---------------- Receive Ports - RX Channel Bonding Ports ----------------
    output          GT2_RXCHANBONDSEQ_OUT,
    input           GT2_RXCHBONDEN_IN,
    input   [2:0]   GT2_RXCHBONDLEVEL_IN,
    input           GT2_RXCHBONDMASTER_IN,
    output  [4:0]   GT2_RXCHBONDO_OUT,
    input           GT2_RXCHBONDSLAVE_IN,
    //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
    output          GT2_RXCHANISALIGNED_OUT,
    output          GT2_RXCHANREALIGN_OUT,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           GT2_GTRXRESET_IN,
    input           GT2_RXPMARESET_IN,
    //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    output  [1:0]   GT2_RXCHARISK_OUT,
    //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
    input   [4:0]   GT2_RXCHBONDI_IN,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          GT2_RXRESETDONE_OUT,
    //------------------- TX Initialization and Reset Ports --------------------
    input           GT2_GTTXRESET_IN,
    input           GT2_TXUSERRDY_IN,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           GT2_TXUSRCLK_IN,
    input           GT2_TXUSRCLK2_IN,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [15:0]  GT2_TXDATA_IN,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          GT2_GTXTXN_OUT,
    output          GT2_GTXTXP_OUT,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          GT2_TXOUTCLK_OUT,
    output          GT2_TXOUTCLKFABRIC_OUT,
    output          GT2_TXOUTCLKPCS_OUT,
    //------------------- Transmit Ports - TX Gearbox Ports --------------------
    input   [1:0]   GT2_TXCHARISK_IN,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    output          GT2_TXRESETDONE_OUT,

    //GT3  (X1Y3)
    //____________________________CHANNEL PORTS________________________________
    //------------------------------- CPLL Ports -------------------------------
    output          GT3_CPLLFBCLKLOST_OUT,
    output          GT3_CPLLLOCK_OUT,
    input           GT3_CPLLLOCKDETCLK_IN,
    input           GT3_CPLLRESET_IN,
    //------------------------ Channel - Clocking Ports ------------------------
    input           GT3_GTREFCLK0_IN,
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   GT3_DRPADDR_IN,
    input           GT3_DRPCLK_IN,
    input   [15:0]  GT3_DRPDI_IN,
    output  [15:0]  GT3_DRPDO_OUT,
    input           GT3_DRPEN_IN,
    output          GT3_DRPRDY_OUT,
    input           GT3_DRPWE_IN,
    //----------------------------- Loopback Ports -----------------------------
    input   [2:0]   GT3_LOOPBACK_IN,
    //------------------- RX Initialization and Reset Ports --------------------
    input           GT3_RXUSERRDY_IN,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          GT3_EYESCANDATAERROR_OUT,
    //----------------------- Receive Ports - CDR Ports ------------------------
    output          GT3_RXCDRLOCK_OUT,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           GT3_RXUSRCLK_IN,
    input           GT3_RXUSRCLK2_IN,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [15:0]  GT3_RXDATA_OUT,
    //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
    output  [1:0]   GT3_RXDISPERR_OUT,
    output  [1:0]   GT3_RXNOTINTABLE_OUT,
    //------------------------- Receive Ports - RX AFE -------------------------
    input           GT3_GTXRXP_IN,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           GT3_GTXRXN_IN,
    //---------------- Receive Ports - RX Channel Bonding Ports ----------------
    output          GT3_RXCHANBONDSEQ_OUT,
    input           GT3_RXCHBONDEN_IN,
    input   [2:0]   GT3_RXCHBONDLEVEL_IN,
    input           GT3_RXCHBONDMASTER_IN,
    output  [4:0]   GT3_RXCHBONDO_OUT,
    input           GT3_RXCHBONDSLAVE_IN,
    //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
    output          GT3_RXCHANISALIGNED_OUT,
    output          GT3_RXCHANREALIGN_OUT,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           GT3_GTRXRESET_IN,
    input           GT3_RXPMARESET_IN,
    //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    output  [1:0]   GT3_RXCHARISK_OUT,
    //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
    input   [4:0]   GT3_RXCHBONDI_IN,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          GT3_RXRESETDONE_OUT,
    //------------------- TX Initialization and Reset Ports --------------------
    input           GT3_GTTXRESET_IN,
    input           GT3_TXUSERRDY_IN,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           GT3_TXUSRCLK_IN,
    input           GT3_TXUSRCLK2_IN,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [15:0]  GT3_TXDATA_IN,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          GT3_GTXTXN_OUT,
    output          GT3_GTXTXP_OUT,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          GT3_TXOUTCLK_OUT,
    output          GT3_TXOUTCLKFABRIC_OUT,
    output          GT3_TXOUTCLKPCS_OUT,
    //------------------- Transmit Ports - TX Gearbox Ports --------------------
    input   [1:0]   GT3_TXCHARISK_IN,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    output          GT3_TXRESETDONE_OUT,

    //GT4  (X1Y8)
    //____________________________CHANNEL PORTS________________________________
    //------------------------------- CPLL Ports -------------------------------
    output          GT4_CPLLFBCLKLOST_OUT,
    output          GT4_CPLLLOCK_OUT,
    input           GT4_CPLLLOCKDETCLK_IN,
    input           GT4_CPLLRESET_IN,
    //------------------------ Channel - Clocking Ports ------------------------
    input           GT4_GTREFCLK0_IN,
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   GT4_DRPADDR_IN,
    input           GT4_DRPCLK_IN,
    input   [15:0]  GT4_DRPDI_IN,
    output  [15:0]  GT4_DRPDO_OUT,
    input           GT4_DRPEN_IN,
    output          GT4_DRPRDY_OUT,
    input           GT4_DRPWE_IN,
    //----------------------------- Loopback Ports -----------------------------
    input   [2:0]   GT4_LOOPBACK_IN,
    //------------------- RX Initialization and Reset Ports --------------------
    input           GT4_RXUSERRDY_IN,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          GT4_EYESCANDATAERROR_OUT,
    //----------------------- Receive Ports - CDR Ports ------------------------
    output          GT4_RXCDRLOCK_OUT,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           GT4_RXUSRCLK_IN,
    input           GT4_RXUSRCLK2_IN,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [15:0]  GT4_RXDATA_OUT,
    //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
    output  [1:0]   GT4_RXDISPERR_OUT,
    output  [1:0]   GT4_RXNOTINTABLE_OUT,
    //------------------------- Receive Ports - RX AFE -------------------------
    input           GT4_GTXRXP_IN,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           GT4_GTXRXN_IN,
    //---------------- Receive Ports - RX Channel Bonding Ports ----------------
    output          GT4_RXCHANBONDSEQ_OUT,
    input           GT4_RXCHBONDEN_IN,
    input   [2:0]   GT4_RXCHBONDLEVEL_IN,
    input           GT4_RXCHBONDMASTER_IN,
    output  [4:0]   GT4_RXCHBONDO_OUT,
    input           GT4_RXCHBONDSLAVE_IN,
    //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
    output          GT4_RXCHANISALIGNED_OUT,
    output          GT4_RXCHANREALIGN_OUT,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           GT4_GTRXRESET_IN,
    input           GT4_RXPMARESET_IN,
    //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    output  [1:0]   GT4_RXCHARISK_OUT,
    //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
    input   [4:0]   GT4_RXCHBONDI_IN,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          GT4_RXRESETDONE_OUT,
    //------------------- TX Initialization and Reset Ports --------------------
    input           GT4_GTTXRESET_IN,
    input           GT4_TXUSERRDY_IN,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           GT4_TXUSRCLK_IN,
    input           GT4_TXUSRCLK2_IN,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [15:0]  GT4_TXDATA_IN,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          GT4_GTXTXN_OUT,
    output          GT4_GTXTXP_OUT,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          GT4_TXOUTCLK_OUT,
    output          GT4_TXOUTCLKFABRIC_OUT,
    output          GT4_TXOUTCLKPCS_OUT,
    //------------------- Transmit Ports - TX Gearbox Ports --------------------
    input   [1:0]   GT4_TXCHARISK_IN,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    output          GT4_TXRESETDONE_OUT,

    //GT5  (X1Y9)
    //____________________________CHANNEL PORTS________________________________
    //------------------------------- CPLL Ports -------------------------------
    output          GT5_CPLLFBCLKLOST_OUT,
    output          GT5_CPLLLOCK_OUT,
    input           GT5_CPLLLOCKDETCLK_IN,
    input           GT5_CPLLRESET_IN,
    //------------------------ Channel - Clocking Ports ------------------------
    input           GT5_GTREFCLK0_IN,
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   GT5_DRPADDR_IN,
    input           GT5_DRPCLK_IN,
    input   [15:0]  GT5_DRPDI_IN,
    output  [15:0]  GT5_DRPDO_OUT,
    input           GT5_DRPEN_IN,
    output          GT5_DRPRDY_OUT,
    input           GT5_DRPWE_IN,
    //----------------------------- Loopback Ports -----------------------------
    input   [2:0]   GT5_LOOPBACK_IN,
    //------------------- RX Initialization and Reset Ports --------------------
    input           GT5_RXUSERRDY_IN,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          GT5_EYESCANDATAERROR_OUT,
    //----------------------- Receive Ports - CDR Ports ------------------------
    output          GT5_RXCDRLOCK_OUT,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           GT5_RXUSRCLK_IN,
    input           GT5_RXUSRCLK2_IN,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [15:0]  GT5_RXDATA_OUT,
    //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
    output  [1:0]   GT5_RXDISPERR_OUT,
    output  [1:0]   GT5_RXNOTINTABLE_OUT,
    //------------------------- Receive Ports - RX AFE -------------------------
    input           GT5_GTXRXP_IN,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           GT5_GTXRXN_IN,
    //---------------- Receive Ports - RX Channel Bonding Ports ----------------
    output          GT5_RXCHANBONDSEQ_OUT,
    input           GT5_RXCHBONDEN_IN,
    input   [2:0]   GT5_RXCHBONDLEVEL_IN,
    input           GT5_RXCHBONDMASTER_IN,
    output  [4:0]   GT5_RXCHBONDO_OUT,
    input           GT5_RXCHBONDSLAVE_IN,
    //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
    output          GT5_RXCHANISALIGNED_OUT,
    output          GT5_RXCHANREALIGN_OUT,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           GT5_GTRXRESET_IN,
    input           GT5_RXPMARESET_IN,
    //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    output  [1:0]   GT5_RXCHARISK_OUT,
    //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
    input   [4:0]   GT5_RXCHBONDI_IN,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          GT5_RXRESETDONE_OUT,
    //------------------- TX Initialization and Reset Ports --------------------
    input           GT5_GTTXRESET_IN,
    input           GT5_TXUSERRDY_IN,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           GT5_TXUSRCLK_IN,
    input           GT5_TXUSRCLK2_IN,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [15:0]  GT5_TXDATA_IN,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          GT5_GTXTXN_OUT,
    output          GT5_GTXTXP_OUT,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          GT5_TXOUTCLK_OUT,
    output          GT5_TXOUTCLKFABRIC_OUT,
    output          GT5_TXOUTCLKPCS_OUT,
    //------------------- Transmit Ports - TX Gearbox Ports --------------------
    input   [1:0]   GT5_TXCHARISK_IN,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    output          GT5_TXRESETDONE_OUT,

    //GT6  (X1Y10)
    //____________________________CHANNEL PORTS________________________________
    //------------------------------- CPLL Ports -------------------------------
    output          GT6_CPLLFBCLKLOST_OUT,
    output          GT6_CPLLLOCK_OUT,
    input           GT6_CPLLLOCKDETCLK_IN,
    input           GT6_CPLLRESET_IN,
    //------------------------ Channel - Clocking Ports ------------------------
    input           GT6_GTREFCLK0_IN,
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   GT6_DRPADDR_IN,
    input           GT6_DRPCLK_IN,
    input   [15:0]  GT6_DRPDI_IN,
    output  [15:0]  GT6_DRPDO_OUT,
    input           GT6_DRPEN_IN,
    output          GT6_DRPRDY_OUT,
    input           GT6_DRPWE_IN,
    //----------------------------- Loopback Ports -----------------------------
    input   [2:0]   GT6_LOOPBACK_IN,
    //------------------- RX Initialization and Reset Ports --------------------
    input           GT6_RXUSERRDY_IN,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          GT6_EYESCANDATAERROR_OUT,
    //----------------------- Receive Ports - CDR Ports ------------------------
    output          GT6_RXCDRLOCK_OUT,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           GT6_RXUSRCLK_IN,
    input           GT6_RXUSRCLK2_IN,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [15:0]  GT6_RXDATA_OUT,
    //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
    output  [1:0]   GT6_RXDISPERR_OUT,
    output  [1:0]   GT6_RXNOTINTABLE_OUT,
    //------------------------- Receive Ports - RX AFE -------------------------
    input           GT6_GTXRXP_IN,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           GT6_GTXRXN_IN,
    //---------------- Receive Ports - RX Channel Bonding Ports ----------------
    output          GT6_RXCHANBONDSEQ_OUT,
    input           GT6_RXCHBONDEN_IN,
    input   [2:0]   GT6_RXCHBONDLEVEL_IN,
    input           GT6_RXCHBONDMASTER_IN,
    output  [4:0]   GT6_RXCHBONDO_OUT,
    input           GT6_RXCHBONDSLAVE_IN,
    //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
    output          GT6_RXCHANISALIGNED_OUT,
    output          GT6_RXCHANREALIGN_OUT,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           GT6_GTRXRESET_IN,
    input           GT6_RXPMARESET_IN,
    //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    output  [1:0]   GT6_RXCHARISK_OUT,
    //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
    input   [4:0]   GT6_RXCHBONDI_IN,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          GT6_RXRESETDONE_OUT,
    //------------------- TX Initialization and Reset Ports --------------------
    input           GT6_GTTXRESET_IN,
    input           GT6_TXUSERRDY_IN,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           GT6_TXUSRCLK_IN,
    input           GT6_TXUSRCLK2_IN,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [15:0]  GT6_TXDATA_IN,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          GT6_GTXTXN_OUT,
    output          GT6_GTXTXP_OUT,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          GT6_TXOUTCLK_OUT,
    output          GT6_TXOUTCLKFABRIC_OUT,
    output          GT6_TXOUTCLKPCS_OUT,
    //------------------- Transmit Ports - TX Gearbox Ports --------------------
    input   [1:0]   GT6_TXCHARISK_IN,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    output          GT6_TXRESETDONE_OUT,

    //GT7  (X1Y11)
    //____________________________CHANNEL PORTS________________________________
    //------------------------------- CPLL Ports -------------------------------
    output          GT7_CPLLFBCLKLOST_OUT,
    output          GT7_CPLLLOCK_OUT,
    input           GT7_CPLLLOCKDETCLK_IN,
    input           GT7_CPLLRESET_IN,
    //------------------------ Channel - Clocking Ports ------------------------
    input           GT7_GTREFCLK0_IN,
    //-------------------------- Channel - DRP Ports  --------------------------
    input   [8:0]   GT7_DRPADDR_IN,
    input           GT7_DRPCLK_IN,
    input   [15:0]  GT7_DRPDI_IN,
    output  [15:0]  GT7_DRPDO_OUT,
    input           GT7_DRPEN_IN,
    output          GT7_DRPRDY_OUT,
    input           GT7_DRPWE_IN,
    //----------------------------- Loopback Ports -----------------------------
    input   [2:0]   GT7_LOOPBACK_IN,
    //------------------- RX Initialization and Reset Ports --------------------
    input           GT7_RXUSERRDY_IN,
    //------------------------ RX Margin Analysis Ports ------------------------
    output          GT7_EYESCANDATAERROR_OUT,
    //----------------------- Receive Ports - CDR Ports ------------------------
    output          GT7_RXCDRLOCK_OUT,
    //---------------- Receive Ports - FPGA RX Interface Ports -----------------
    input           GT7_RXUSRCLK_IN,
    input           GT7_RXUSRCLK2_IN,
    //---------------- Receive Ports - FPGA RX interface Ports -----------------
    output  [15:0]  GT7_RXDATA_OUT,
    //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
    output  [1:0]   GT7_RXDISPERR_OUT,
    output  [1:0]   GT7_RXNOTINTABLE_OUT,
    //------------------------- Receive Ports - RX AFE -------------------------
    input           GT7_GTXRXP_IN,
    //---------------------- Receive Ports - RX AFE Ports ----------------------
    input           GT7_GTXRXN_IN,
    //---------------- Receive Ports - RX Channel Bonding Ports ----------------
    output          GT7_RXCHANBONDSEQ_OUT,
    input           GT7_RXCHBONDEN_IN,
    input   [2:0]   GT7_RXCHBONDLEVEL_IN,
    input           GT7_RXCHBONDMASTER_IN,
    output  [4:0]   GT7_RXCHBONDO_OUT,
    input           GT7_RXCHBONDSLAVE_IN,
    //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
    output          GT7_RXCHANISALIGNED_OUT,
    output          GT7_RXCHANREALIGN_OUT,
    //----------- Receive Ports - RX Initialization and Reset Ports ------------
    input           GT7_GTRXRESET_IN,
    input           GT7_RXPMARESET_IN,
    //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
    output  [1:0]   GT7_RXCHARISK_OUT,
    //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
    input   [4:0]   GT7_RXCHBONDI_IN,
    //------------ Receive Ports -RX Initialization and Reset Ports ------------
    output          GT7_RXRESETDONE_OUT,
    //------------------- TX Initialization and Reset Ports --------------------
    input           GT7_GTTXRESET_IN,
    input           GT7_TXUSERRDY_IN,
    //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
    input           GT7_TXUSRCLK_IN,
    input           GT7_TXUSRCLK2_IN,
    //---------------- Transmit Ports - TX Data Path interface -----------------
    input   [15:0]  GT7_TXDATA_IN,
    //-------------- Transmit Ports - TX Driver and OOB signaling --------------
    output          GT7_GTXTXN_OUT,
    output          GT7_GTXTXP_OUT,
    //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    output          GT7_TXOUTCLK_OUT,
    output          GT7_TXOUTCLKFABRIC_OUT,
    output          GT7_TXOUTCLKPCS_OUT,
    //------------------- Transmit Ports - TX Gearbox Ports --------------------
    input   [1:0]   GT7_TXCHARISK_IN,
    //----------- Transmit Ports - TX Initialization and Reset Ports -----------
    output          GT7_TXRESETDONE_OUT,


    //____________________________COMMON PORTS________________________________
    //-------------------- Common Block  - Ref Clock Ports ---------------------
    input           GT0_GTREFCLK0_COMMON_IN,
    //----------------------- Common Block - QPLL Ports ------------------------
    output          GT0_QPLLLOCK_OUT,
    input           GT0_QPLLLOCKDETCLK_IN,
    input           GT0_QPLLRESET_IN,

    //____________________________COMMON PORTS________________________________
    //-------------------- Common Block  - Ref Clock Ports ---------------------
    input           GT1_GTREFCLK0_COMMON_IN,
    //----------------------- Common Block - QPLL Ports ------------------------
    output          GT1_QPLLLOCK_OUT,
    input           GT1_QPLLLOCKDETCLK_IN,
    input           GT1_QPLLRESET_IN


);



//***********************************Parameter Declarations********************

    //Typical CDRLOCK Time is 50,000UI, as per DS183
    parameter RX_CDRLOCK_TIME      = (EXAMPLE_SIMULATION == 1) ? 1000 : 50000/3.125;

       
    integer   WAIT_TIME_CDRLOCK    = RX_CDRLOCK_TIME / STABLE_CLOCK_PERIOD;      

//-------------------------- GT Wrapper Wires ------------------------------
    wire           gt0_cpllreset_i;
    wire           gt0_cpllreset_t;
    wire           gt0_cpllrefclklost_i;
    wire           gt0_cplllock_i;
    wire           gt0_txresetdone_i;
    wire           gt0_rxresetdone_i;
    wire           gt0_gttxreset_i;
    wire           gt0_gttxreset_t;
    wire           gt0_gtrxreset_i;
    wire           gt0_gtrxreset_t;
    wire           gt0_rxdfelpmreset_i;
    wire           gt0_txuserrdy_i;
    wire           gt0_txuserrdy_t;
    wire           gt0_rxuserrdy_i;
    wire           gt0_rxuserrdy_t;

    wire           gt0_rxdfeagchold_i;
    wire           gt0_rxdfelfhold_i;
    wire           gt0_rxlpmlfhold_i;
    wire           gt0_rxlpmhfhold_i;


    wire           gt1_cpllreset_i;
    wire           gt1_cpllreset_t;
    wire           gt1_cpllrefclklost_i;
    wire           gt1_cplllock_i;
    wire           gt1_txresetdone_i;
    wire           gt1_rxresetdone_i;
    wire           gt1_gttxreset_i;
    wire           gt1_gttxreset_t;
    wire           gt1_gtrxreset_i;
    wire           gt1_gtrxreset_t;
    wire           gt1_rxdfelpmreset_i;
    wire           gt1_txuserrdy_i;
    wire           gt1_txuserrdy_t;
    wire           gt1_rxuserrdy_i;
    wire           gt1_rxuserrdy_t;

    wire           gt1_rxdfeagchold_i;
    wire           gt1_rxdfelfhold_i;
    wire           gt1_rxlpmlfhold_i;
    wire           gt1_rxlpmhfhold_i;


    wire           gt2_cpllreset_i;
    wire           gt2_cpllreset_t;
    wire           gt2_cpllrefclklost_i;
    wire           gt2_cplllock_i;
    wire           gt2_txresetdone_i;
    wire           gt2_rxresetdone_i;
    wire           gt2_gttxreset_i;
    wire           gt2_gttxreset_t;
    wire           gt2_gtrxreset_i;
    wire           gt2_gtrxreset_t;
    wire           gt2_rxdfelpmreset_i;
    wire           gt2_txuserrdy_i;
    wire           gt2_txuserrdy_t;
    wire           gt2_rxuserrdy_i;
    wire           gt2_rxuserrdy_t;

    wire           gt2_rxdfeagchold_i;
    wire           gt2_rxdfelfhold_i;
    wire           gt2_rxlpmlfhold_i;
    wire           gt2_rxlpmhfhold_i;


    wire           gt3_cpllreset_i;
    wire           gt3_cpllreset_t;
    wire           gt3_cpllrefclklost_i;
    wire           gt3_cplllock_i;
    wire           gt3_txresetdone_i;
    wire           gt3_rxresetdone_i;
    wire           gt3_gttxreset_i;
    wire           gt3_gttxreset_t;
    wire           gt3_gtrxreset_i;
    wire           gt3_gtrxreset_t;
    wire           gt3_rxdfelpmreset_i;
    wire           gt3_txuserrdy_i;
    wire           gt3_txuserrdy_t;
    wire           gt3_rxuserrdy_i;
    wire           gt3_rxuserrdy_t;

    wire           gt3_rxdfeagchold_i;
    wire           gt3_rxdfelfhold_i;
    wire           gt3_rxlpmlfhold_i;
    wire           gt3_rxlpmhfhold_i;


    wire           gt4_cpllreset_i;
    wire           gt4_cpllreset_t;
    wire           gt4_cpllrefclklost_i;
    wire           gt4_cplllock_i;
    wire           gt4_txresetdone_i;
    wire           gt4_rxresetdone_i;
    wire           gt4_gttxreset_i;
    wire           gt4_gttxreset_t;
    wire           gt4_gtrxreset_i;
    wire           gt4_gtrxreset_t;
    wire           gt4_rxdfelpmreset_i;
    wire           gt4_txuserrdy_i;
    wire           gt4_txuserrdy_t;
    wire           gt4_rxuserrdy_i;
    wire           gt4_rxuserrdy_t;

    wire           gt4_rxdfeagchold_i;
    wire           gt4_rxdfelfhold_i;
    wire           gt4_rxlpmlfhold_i;
    wire           gt4_rxlpmhfhold_i;


    wire           gt5_cpllreset_i;
    wire           gt5_cpllreset_t;
    wire           gt5_cpllrefclklost_i;
    wire           gt5_cplllock_i;
    wire           gt5_txresetdone_i;
    wire           gt5_rxresetdone_i;
    wire           gt5_gttxreset_i;
    wire           gt5_gttxreset_t;
    wire           gt5_gtrxreset_i;
    wire           gt5_gtrxreset_t;
    wire           gt5_rxdfelpmreset_i;
    wire           gt5_txuserrdy_i;
    wire           gt5_txuserrdy_t;
    wire           gt5_rxuserrdy_i;
    wire           gt5_rxuserrdy_t;

    wire           gt5_rxdfeagchold_i;
    wire           gt5_rxdfelfhold_i;
    wire           gt5_rxlpmlfhold_i;
    wire           gt5_rxlpmhfhold_i;


    wire           gt6_cpllreset_i;
    wire           gt6_cpllreset_t;
    wire           gt6_cpllrefclklost_i;
    wire           gt6_cplllock_i;
    wire           gt6_txresetdone_i;
    wire           gt6_rxresetdone_i;
    wire           gt6_gttxreset_i;
    wire           gt6_gttxreset_t;
    wire           gt6_gtrxreset_i;
    wire           gt6_gtrxreset_t;
    wire           gt6_rxdfelpmreset_i;
    wire           gt6_txuserrdy_i;
    wire           gt6_txuserrdy_t;
    wire           gt6_rxuserrdy_i;
    wire           gt6_rxuserrdy_t;

    wire           gt6_rxdfeagchold_i;
    wire           gt6_rxdfelfhold_i;
    wire           gt6_rxlpmlfhold_i;
    wire           gt6_rxlpmhfhold_i;


    wire           gt7_cpllreset_i;
    wire           gt7_cpllreset_t;
    wire           gt7_cpllrefclklost_i;
    wire           gt7_cplllock_i;
    wire           gt7_txresetdone_i;
    wire           gt7_rxresetdone_i;
    wire           gt7_gttxreset_i;
    wire           gt7_gttxreset_t;
    wire           gt7_gtrxreset_i;
    wire           gt7_gtrxreset_t;
    wire           gt7_rxdfelpmreset_i;
    wire           gt7_txuserrdy_i;
    wire           gt7_txuserrdy_t;
    wire           gt7_rxuserrdy_i;
    wire           gt7_rxuserrdy_t;

    wire           gt7_rxdfeagchold_i;
    wire           gt7_rxdfelfhold_i;
    wire           gt7_rxlpmlfhold_i;
    wire           gt7_rxlpmhfhold_i;



    wire           gt0_qpllreset_i;
    wire           gt0_qpllreset_t;
    wire           gt0_qpllrefclklost_i;
    wire           gt0_qplllock_i;
    wire           gt1_qpllreset_i;
    wire           gt1_qpllreset_t;
    wire           gt1_qpllrefclklost_i;
    wire           gt1_qplllock_i;


//------------------------------- Global Signals -----------------------------
    wire           tied_to_ground_i;
    wire           tied_to_vcc_i;

    wire           gt0_rxoutclk_i;
    wire           gt0_recclk_stable_i;

    wire           gt1_rxoutclk_i;
    wire           gt1_recclk_stable_i;

    wire           gt2_rxoutclk_i;
    wire           gt2_recclk_stable_i;

    wire           gt3_rxoutclk_i;
    wire           gt3_recclk_stable_i;

    wire           gt4_rxoutclk_i;
    wire           gt4_recclk_stable_i;

    wire           gt5_rxoutclk_i;
    wire           gt5_recclk_stable_i;

    wire           gt6_rxoutclk_i;
    wire           gt6_recclk_stable_i;

    wire           gt7_rxoutclk_i;
    wire           gt7_recclk_stable_i;







    integer  rx_cdrlock_counter= 0;
    reg              rx_cdrlocked;


 


//**************************** Main Body of Code *******************************
    //  Static signal Assigments
    assign  tied_to_ground_i                     =  1'b0;
    assign  tied_to_vcc_i                        =  1'b1;

//    ----------------------------- The GT Wrapper -----------------------------
    
    // Use the instantiation template in the example directory to add the GT wrapper to your design.
    // In this example, the wrapper is wired up for basic operation with a frame generator and frame 
    // checker. The GTs will reset, then attempt to align and transmit data. If channel bonding is 
    // enabled, bonding should occur after alignment.


    serdes_coe #
    (
        .WRAPPER_SIM_GTRESET_SPEEDUP    (EXAMPLE_SIM_GTRESET_SPEEDUP)
    )
    serdes_coe_i
    (
  
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT0  (X1Y0)

        //------------------------------- CPLL Ports -------------------------------
        .GT0_CPLLFBCLKLOST_OUT          (GT0_CPLLFBCLKLOST_OUT),
        .GT0_CPLLLOCK_OUT               (gt0_cplllock_i),
        .GT0_CPLLLOCKDETCLK_IN          (GT0_CPLLLOCKDETCLK_IN),
        .GT0_CPLLREFCLKLOST_OUT         (gt0_cpllrefclklost_i),
        .GT0_CPLLRESET_IN               (gt0_cpllreset_i),
        //------------------------ Channel - Clocking Ports ------------------------
        .GT0_GTREFCLK0_IN               (GT0_GTREFCLK0_IN),
        //-------------------------- Channel - DRP Ports  --------------------------
        .GT0_DRPADDR_IN                 (GT0_DRPADDR_IN),
        .GT0_DRPCLK_IN                  (GT0_DRPCLK_IN),
        .GT0_DRPDI_IN                   (GT0_DRPDI_IN),
        .GT0_DRPDO_OUT                  (GT0_DRPDO_OUT),
        .GT0_DRPEN_IN                   (GT0_DRPEN_IN),
        .GT0_DRPRDY_OUT                 (GT0_DRPRDY_OUT),
        .GT0_DRPWE_IN                   (GT0_DRPWE_IN),
        //----------------------------- Loopback Ports -----------------------------
        .GT0_LOOPBACK_IN                (GT0_LOOPBACK_IN),
        //------------------- RX Initialization and Reset Ports --------------------
        .GT0_RXUSERRDY_IN               (gt0_rxuserrdy_i),
        //------------------------ RX Margin Analysis Ports ------------------------
        .GT0_EYESCANDATAERROR_OUT       (GT0_EYESCANDATAERROR_OUT),
        //----------------------- Receive Ports - CDR Ports ------------------------
        .GT0_RXCDRLOCK_OUT              (GT0_RXCDRLOCK_OUT),
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .GT0_RXUSRCLK_IN                (GT0_RXUSRCLK_IN),
        .GT0_RXUSRCLK2_IN               (GT0_RXUSRCLK2_IN),
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .GT0_RXDATA_OUT                 (GT0_RXDATA_OUT),
        //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
        .GT0_RXDISPERR_OUT              (GT0_RXDISPERR_OUT),
        .GT0_RXNOTINTABLE_OUT           (GT0_RXNOTINTABLE_OUT),
        //------------------------- Receive Ports - RX AFE -------------------------
        .GT0_GTXRXP_IN                  (GT0_GTXRXP_IN),
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .GT0_GTXRXN_IN                  (GT0_GTXRXN_IN),
        //---------------- Receive Ports - RX Channel Bonding Ports ----------------
        .GT0_RXCHANBONDSEQ_OUT          (GT0_RXCHANBONDSEQ_OUT),
        .GT0_RXCHBONDEN_IN              (GT0_RXCHBONDEN_IN),
        .GT0_RXCHBONDLEVEL_IN           (GT0_RXCHBONDLEVEL_IN),
        .GT0_RXCHBONDMASTER_IN          (GT0_RXCHBONDMASTER_IN),
        .GT0_RXCHBONDO_OUT              (GT0_RXCHBONDO_OUT),
        .GT0_RXCHBONDSLAVE_IN           (GT0_RXCHBONDSLAVE_IN),
        //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
        .GT0_RXCHANISALIGNED_OUT        (GT0_RXCHANISALIGNED_OUT),
        .GT0_RXCHANREALIGN_OUT          (GT0_RXCHANREALIGN_OUT),
        //------------------ Receive Ports - RX Equailizer Ports -------------------
        .GT0_RXLPMHFHOLD_IN             (gt0_rxlpmhfhold_i),
        .GT0_RXLPMLFHOLD_IN             (gt0_rxlpmlfhold_i),
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .GT0_RXOUTCLK_OUT               (gt0_rxoutclk_i),
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .GT0_GTRXRESET_IN               (gt0_gtrxreset_i),
        .GT0_RXPMARESET_IN              (GT0_RXPMARESET_IN),
        //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        .GT0_RXCHARISK_OUT              (GT0_RXCHARISK_OUT),
        //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
        .GT0_RXCHBONDI_IN               (GT0_RXCHBONDI_IN),
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .GT0_RXRESETDONE_OUT            (gt0_rxresetdone_i),
        //------------------- TX Initialization and Reset Ports --------------------
        .GT0_GTTXRESET_IN               (gt0_gttxreset_i),
        .GT0_TXUSERRDY_IN               (gt0_txuserrdy_i),
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .GT0_TXUSRCLK_IN                (GT0_TXUSRCLK_IN),
        .GT0_TXUSRCLK2_IN               (GT0_TXUSRCLK2_IN),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .GT0_TXDATA_IN                  (GT0_TXDATA_IN),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .GT0_GTXTXN_OUT                 (GT0_GTXTXN_OUT),
        .GT0_GTXTXP_OUT                 (GT0_GTXTXP_OUT),
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .GT0_TXOUTCLK_OUT               (GT0_TXOUTCLK_OUT),
        .GT0_TXOUTCLKFABRIC_OUT         (GT0_TXOUTCLKFABRIC_OUT),
        .GT0_TXOUTCLKPCS_OUT            (GT0_TXOUTCLKPCS_OUT),
        //------------------- Transmit Ports - TX Gearbox Ports --------------------
        .GT0_TXCHARISK_IN               (GT0_TXCHARISK_IN),
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .GT0_TXRESETDONE_OUT            (gt0_txresetdone_i),


  
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT1  (X1Y1)

        //------------------------------- CPLL Ports -------------------------------
        .GT1_CPLLFBCLKLOST_OUT          (GT1_CPLLFBCLKLOST_OUT),
        .GT1_CPLLLOCK_OUT               (gt1_cplllock_i),
        .GT1_CPLLLOCKDETCLK_IN          (GT1_CPLLLOCKDETCLK_IN),
        .GT1_CPLLREFCLKLOST_OUT         (gt1_cpllrefclklost_i),
        .GT1_CPLLRESET_IN               (gt1_cpllreset_i),
        //------------------------ Channel - Clocking Ports ------------------------
        .GT1_GTREFCLK0_IN               (GT1_GTREFCLK0_IN),
        //-------------------------- Channel - DRP Ports  --------------------------
        .GT1_DRPADDR_IN                 (GT1_DRPADDR_IN),
        .GT1_DRPCLK_IN                  (GT1_DRPCLK_IN),
        .GT1_DRPDI_IN                   (GT1_DRPDI_IN),
        .GT1_DRPDO_OUT                  (GT1_DRPDO_OUT),
        .GT1_DRPEN_IN                   (GT1_DRPEN_IN),
        .GT1_DRPRDY_OUT                 (GT1_DRPRDY_OUT),
        .GT1_DRPWE_IN                   (GT1_DRPWE_IN),
        //----------------------------- Loopback Ports -----------------------------
        .GT1_LOOPBACK_IN                (GT1_LOOPBACK_IN),
        //------------------- RX Initialization and Reset Ports --------------------
        .GT1_RXUSERRDY_IN               (gt1_rxuserrdy_i),
        //------------------------ RX Margin Analysis Ports ------------------------
        .GT1_EYESCANDATAERROR_OUT       (GT1_EYESCANDATAERROR_OUT),
        //----------------------- Receive Ports - CDR Ports ------------------------
        .GT1_RXCDRLOCK_OUT              (GT1_RXCDRLOCK_OUT),
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .GT1_RXUSRCLK_IN                (GT1_RXUSRCLK_IN),
        .GT1_RXUSRCLK2_IN               (GT1_RXUSRCLK2_IN),
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .GT1_RXDATA_OUT                 (GT1_RXDATA_OUT),
        //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
        .GT1_RXDISPERR_OUT              (GT1_RXDISPERR_OUT),
        .GT1_RXNOTINTABLE_OUT           (GT1_RXNOTINTABLE_OUT),
        //------------------------- Receive Ports - RX AFE -------------------------
        .GT1_GTXRXP_IN                  (GT1_GTXRXP_IN),
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .GT1_GTXRXN_IN                  (GT1_GTXRXN_IN),
        //---------------- Receive Ports - RX Channel Bonding Ports ----------------
        .GT1_RXCHANBONDSEQ_OUT          (GT1_RXCHANBONDSEQ_OUT),
        .GT1_RXCHBONDEN_IN              (GT1_RXCHBONDEN_IN),
        .GT1_RXCHBONDLEVEL_IN           (GT1_RXCHBONDLEVEL_IN),
        .GT1_RXCHBONDMASTER_IN          (GT1_RXCHBONDMASTER_IN),
        .GT1_RXCHBONDO_OUT              (GT1_RXCHBONDO_OUT),
        .GT1_RXCHBONDSLAVE_IN           (GT1_RXCHBONDSLAVE_IN),
        //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
        .GT1_RXCHANISALIGNED_OUT        (GT1_RXCHANISALIGNED_OUT),
        .GT1_RXCHANREALIGN_OUT          (GT1_RXCHANREALIGN_OUT),
        //------------------ Receive Ports - RX Equailizer Ports -------------------
        .GT1_RXLPMHFHOLD_IN             (gt1_rxlpmhfhold_i),
        .GT1_RXLPMLFHOLD_IN             (gt1_rxlpmlfhold_i),
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .GT1_RXOUTCLK_OUT               (gt1_rxoutclk_i),
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .GT1_GTRXRESET_IN               (gt1_gtrxreset_i),
        .GT1_RXPMARESET_IN              (GT1_RXPMARESET_IN),
        //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        .GT1_RXCHARISK_OUT              (GT1_RXCHARISK_OUT),
        //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
        .GT1_RXCHBONDI_IN               (GT1_RXCHBONDI_IN),
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .GT1_RXRESETDONE_OUT            (gt1_rxresetdone_i),
        //------------------- TX Initialization and Reset Ports --------------------
        .GT1_GTTXRESET_IN               (gt1_gttxreset_i),
        .GT1_TXUSERRDY_IN               (gt1_txuserrdy_i),
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .GT1_TXUSRCLK_IN                (GT1_TXUSRCLK_IN),
        .GT1_TXUSRCLK2_IN               (GT1_TXUSRCLK2_IN),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .GT1_TXDATA_IN                  (GT1_TXDATA_IN),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .GT1_GTXTXN_OUT                 (GT1_GTXTXN_OUT),
        .GT1_GTXTXP_OUT                 (GT1_GTXTXP_OUT),
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .GT1_TXOUTCLK_OUT               (GT1_TXOUTCLK_OUT),
        .GT1_TXOUTCLKFABRIC_OUT         (GT1_TXOUTCLKFABRIC_OUT),
        .GT1_TXOUTCLKPCS_OUT            (GT1_TXOUTCLKPCS_OUT),
        //------------------- Transmit Ports - TX Gearbox Ports --------------------
        .GT1_TXCHARISK_IN               (GT1_TXCHARISK_IN),
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .GT1_TXRESETDONE_OUT            (gt1_txresetdone_i),


  
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT2  (X1Y2)

        //------------------------------- CPLL Ports -------------------------------
        .GT2_CPLLFBCLKLOST_OUT          (GT2_CPLLFBCLKLOST_OUT),
        .GT2_CPLLLOCK_OUT               (gt2_cplllock_i),
        .GT2_CPLLLOCKDETCLK_IN          (GT2_CPLLLOCKDETCLK_IN),
        .GT2_CPLLREFCLKLOST_OUT         (gt2_cpllrefclklost_i),
        .GT2_CPLLRESET_IN               (gt2_cpllreset_i),
        //------------------------ Channel - Clocking Ports ------------------------
        .GT2_GTREFCLK0_IN               (GT2_GTREFCLK0_IN),
        //-------------------------- Channel - DRP Ports  --------------------------
        .GT2_DRPADDR_IN                 (GT2_DRPADDR_IN),
        .GT2_DRPCLK_IN                  (GT2_DRPCLK_IN),
        .GT2_DRPDI_IN                   (GT2_DRPDI_IN),
        .GT2_DRPDO_OUT                  (GT2_DRPDO_OUT),
        .GT2_DRPEN_IN                   (GT2_DRPEN_IN),
        .GT2_DRPRDY_OUT                 (GT2_DRPRDY_OUT),
        .GT2_DRPWE_IN                   (GT2_DRPWE_IN),
        //----------------------------- Loopback Ports -----------------------------
        .GT2_LOOPBACK_IN                (GT2_LOOPBACK_IN),
        //------------------- RX Initialization and Reset Ports --------------------
        .GT2_RXUSERRDY_IN               (gt2_rxuserrdy_i),
        //------------------------ RX Margin Analysis Ports ------------------------
        .GT2_EYESCANDATAERROR_OUT       (GT2_EYESCANDATAERROR_OUT),
        //----------------------- Receive Ports - CDR Ports ------------------------
        .GT2_RXCDRLOCK_OUT              (GT2_RXCDRLOCK_OUT),
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .GT2_RXUSRCLK_IN                (GT2_RXUSRCLK_IN),
        .GT2_RXUSRCLK2_IN               (GT2_RXUSRCLK2_IN),
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .GT2_RXDATA_OUT                 (GT2_RXDATA_OUT),
        //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
        .GT2_RXDISPERR_OUT              (GT2_RXDISPERR_OUT),
        .GT2_RXNOTINTABLE_OUT           (GT2_RXNOTINTABLE_OUT),
        //------------------------- Receive Ports - RX AFE -------------------------
        .GT2_GTXRXP_IN                  (GT2_GTXRXP_IN),
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .GT2_GTXRXN_IN                  (GT2_GTXRXN_IN),
        //---------------- Receive Ports - RX Channel Bonding Ports ----------------
        .GT2_RXCHANBONDSEQ_OUT          (GT2_RXCHANBONDSEQ_OUT),
        .GT2_RXCHBONDEN_IN              (GT2_RXCHBONDEN_IN),
        .GT2_RXCHBONDLEVEL_IN           (GT2_RXCHBONDLEVEL_IN),
        .GT2_RXCHBONDMASTER_IN          (GT2_RXCHBONDMASTER_IN),
        .GT2_RXCHBONDO_OUT              (GT2_RXCHBONDO_OUT),
        .GT2_RXCHBONDSLAVE_IN           (GT2_RXCHBONDSLAVE_IN),
        //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
        .GT2_RXCHANISALIGNED_OUT        (GT2_RXCHANISALIGNED_OUT),
        .GT2_RXCHANREALIGN_OUT          (GT2_RXCHANREALIGN_OUT),
        //------------------ Receive Ports - RX Equailizer Ports -------------------
        .GT2_RXLPMHFHOLD_IN             (gt2_rxlpmhfhold_i),
        .GT2_RXLPMLFHOLD_IN             (gt2_rxlpmlfhold_i),
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .GT2_RXOUTCLK_OUT               (gt2_rxoutclk_i),
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .GT2_GTRXRESET_IN               (gt2_gtrxreset_i),
        .GT2_RXPMARESET_IN              (GT2_RXPMARESET_IN),
        //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        .GT2_RXCHARISK_OUT              (GT2_RXCHARISK_OUT),
        //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
        .GT2_RXCHBONDI_IN               (GT2_RXCHBONDI_IN),
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .GT2_RXRESETDONE_OUT            (gt2_rxresetdone_i),
        //------------------- TX Initialization and Reset Ports --------------------
        .GT2_GTTXRESET_IN               (gt2_gttxreset_i),
        .GT2_TXUSERRDY_IN               (gt2_txuserrdy_i),
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .GT2_TXUSRCLK_IN                (GT2_TXUSRCLK_IN),
        .GT2_TXUSRCLK2_IN               (GT2_TXUSRCLK2_IN),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .GT2_TXDATA_IN                  (GT2_TXDATA_IN),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .GT2_GTXTXN_OUT                 (GT2_GTXTXN_OUT),
        .GT2_GTXTXP_OUT                 (GT2_GTXTXP_OUT),
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .GT2_TXOUTCLK_OUT               (GT2_TXOUTCLK_OUT),
        .GT2_TXOUTCLKFABRIC_OUT         (GT2_TXOUTCLKFABRIC_OUT),
        .GT2_TXOUTCLKPCS_OUT            (GT2_TXOUTCLKPCS_OUT),
        //------------------- Transmit Ports - TX Gearbox Ports --------------------
        .GT2_TXCHARISK_IN               (GT2_TXCHARISK_IN),
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .GT2_TXRESETDONE_OUT            (gt2_txresetdone_i),


  
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT3  (X1Y3)

        //------------------------------- CPLL Ports -------------------------------
        .GT3_CPLLFBCLKLOST_OUT          (GT3_CPLLFBCLKLOST_OUT),
        .GT3_CPLLLOCK_OUT               (gt3_cplllock_i),
        .GT3_CPLLLOCKDETCLK_IN          (GT3_CPLLLOCKDETCLK_IN),
        .GT3_CPLLREFCLKLOST_OUT         (gt3_cpllrefclklost_i),
        .GT3_CPLLRESET_IN               (gt3_cpllreset_i),
        //------------------------ Channel - Clocking Ports ------------------------
        .GT3_GTREFCLK0_IN               (GT3_GTREFCLK0_IN),
        //-------------------------- Channel - DRP Ports  --------------------------
        .GT3_DRPADDR_IN                 (GT3_DRPADDR_IN),
        .GT3_DRPCLK_IN                  (GT3_DRPCLK_IN),
        .GT3_DRPDI_IN                   (GT3_DRPDI_IN),
        .GT3_DRPDO_OUT                  (GT3_DRPDO_OUT),
        .GT3_DRPEN_IN                   (GT3_DRPEN_IN),
        .GT3_DRPRDY_OUT                 (GT3_DRPRDY_OUT),
        .GT3_DRPWE_IN                   (GT3_DRPWE_IN),
        //----------------------------- Loopback Ports -----------------------------
        .GT3_LOOPBACK_IN                (GT3_LOOPBACK_IN),
        //------------------- RX Initialization and Reset Ports --------------------
        .GT3_RXUSERRDY_IN               (gt3_rxuserrdy_i),
        //------------------------ RX Margin Analysis Ports ------------------------
        .GT3_EYESCANDATAERROR_OUT       (GT3_EYESCANDATAERROR_OUT),
        //----------------------- Receive Ports - CDR Ports ------------------------
        .GT3_RXCDRLOCK_OUT              (GT3_RXCDRLOCK_OUT),
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .GT3_RXUSRCLK_IN                (GT3_RXUSRCLK_IN),
        .GT3_RXUSRCLK2_IN               (GT3_RXUSRCLK2_IN),
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .GT3_RXDATA_OUT                 (GT3_RXDATA_OUT),
        //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
        .GT3_RXDISPERR_OUT              (GT3_RXDISPERR_OUT),
        .GT3_RXNOTINTABLE_OUT           (GT3_RXNOTINTABLE_OUT),
        //------------------------- Receive Ports - RX AFE -------------------------
        .GT3_GTXRXP_IN                  (GT3_GTXRXP_IN),
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .GT3_GTXRXN_IN                  (GT3_GTXRXN_IN),
        //---------------- Receive Ports - RX Channel Bonding Ports ----------------
        .GT3_RXCHANBONDSEQ_OUT          (GT3_RXCHANBONDSEQ_OUT),
        .GT3_RXCHBONDEN_IN              (GT3_RXCHBONDEN_IN),
        .GT3_RXCHBONDLEVEL_IN           (GT3_RXCHBONDLEVEL_IN),
        .GT3_RXCHBONDMASTER_IN          (GT3_RXCHBONDMASTER_IN),
        .GT3_RXCHBONDO_OUT              (GT3_RXCHBONDO_OUT),
        .GT3_RXCHBONDSLAVE_IN           (GT3_RXCHBONDSLAVE_IN),
        //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
        .GT3_RXCHANISALIGNED_OUT        (GT3_RXCHANISALIGNED_OUT),
        .GT3_RXCHANREALIGN_OUT          (GT3_RXCHANREALIGN_OUT),
        //------------------ Receive Ports - RX Equailizer Ports -------------------
        .GT3_RXLPMHFHOLD_IN             (gt3_rxlpmhfhold_i),
        .GT3_RXLPMLFHOLD_IN             (gt3_rxlpmlfhold_i),
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .GT3_RXOUTCLK_OUT               (gt3_rxoutclk_i),
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .GT3_GTRXRESET_IN               (gt3_gtrxreset_i),
        .GT3_RXPMARESET_IN              (GT3_RXPMARESET_IN),
        //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        .GT3_RXCHARISK_OUT              (GT3_RXCHARISK_OUT),
        //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
        .GT3_RXCHBONDI_IN               (GT3_RXCHBONDI_IN),
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .GT3_RXRESETDONE_OUT            (gt3_rxresetdone_i),
        //------------------- TX Initialization and Reset Ports --------------------
        .GT3_GTTXRESET_IN               (gt3_gttxreset_i),
        .GT3_TXUSERRDY_IN               (gt3_txuserrdy_i),
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .GT3_TXUSRCLK_IN                (GT3_TXUSRCLK_IN),
        .GT3_TXUSRCLK2_IN               (GT3_TXUSRCLK2_IN),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .GT3_TXDATA_IN                  (GT3_TXDATA_IN),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .GT3_GTXTXN_OUT                 (GT3_GTXTXN_OUT),
        .GT3_GTXTXP_OUT                 (GT3_GTXTXP_OUT),
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .GT3_TXOUTCLK_OUT               (GT3_TXOUTCLK_OUT),
        .GT3_TXOUTCLKFABRIC_OUT         (GT3_TXOUTCLKFABRIC_OUT),
        .GT3_TXOUTCLKPCS_OUT            (GT3_TXOUTCLKPCS_OUT),
        //------------------- Transmit Ports - TX Gearbox Ports --------------------
        .GT3_TXCHARISK_IN               (GT3_TXCHARISK_IN),
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .GT3_TXRESETDONE_OUT            (gt3_txresetdone_i),


  
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT4  (X1Y8)

        //------------------------------- CPLL Ports -------------------------------
        .GT4_CPLLFBCLKLOST_OUT          (GT4_CPLLFBCLKLOST_OUT),
        .GT4_CPLLLOCK_OUT               (gt4_cplllock_i),
        .GT4_CPLLLOCKDETCLK_IN          (GT4_CPLLLOCKDETCLK_IN),
        .GT4_CPLLREFCLKLOST_OUT         (gt4_cpllrefclklost_i),
        .GT4_CPLLRESET_IN               (gt4_cpllreset_i),
        //------------------------ Channel - Clocking Ports ------------------------
        .GT4_GTREFCLK0_IN               (GT4_GTREFCLK0_IN),
        //-------------------------- Channel - DRP Ports  --------------------------
        .GT4_DRPADDR_IN                 (GT4_DRPADDR_IN),
        .GT4_DRPCLK_IN                  (GT4_DRPCLK_IN),
        .GT4_DRPDI_IN                   (GT4_DRPDI_IN),
        .GT4_DRPDO_OUT                  (GT4_DRPDO_OUT),
        .GT4_DRPEN_IN                   (GT4_DRPEN_IN),
        .GT4_DRPRDY_OUT                 (GT4_DRPRDY_OUT),
        .GT4_DRPWE_IN                   (GT4_DRPWE_IN),
        //----------------------------- Loopback Ports -----------------------------
        .GT4_LOOPBACK_IN                (GT4_LOOPBACK_IN),
        //------------------- RX Initialization and Reset Ports --------------------
        .GT4_RXUSERRDY_IN               (gt4_rxuserrdy_i),
        //------------------------ RX Margin Analysis Ports ------------------------
        .GT4_EYESCANDATAERROR_OUT       (GT4_EYESCANDATAERROR_OUT),
        //----------------------- Receive Ports - CDR Ports ------------------------
        .GT4_RXCDRLOCK_OUT              (GT4_RXCDRLOCK_OUT),
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .GT4_RXUSRCLK_IN                (GT4_RXUSRCLK_IN),
        .GT4_RXUSRCLK2_IN               (GT4_RXUSRCLK2_IN),
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .GT4_RXDATA_OUT                 (GT4_RXDATA_OUT),
        //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
        .GT4_RXDISPERR_OUT              (GT4_RXDISPERR_OUT),
        .GT4_RXNOTINTABLE_OUT           (GT4_RXNOTINTABLE_OUT),
        //------------------------- Receive Ports - RX AFE -------------------------
        .GT4_GTXRXP_IN                  (GT4_GTXRXP_IN),
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .GT4_GTXRXN_IN                  (GT4_GTXRXN_IN),
        //---------------- Receive Ports - RX Channel Bonding Ports ----------------
        .GT4_RXCHANBONDSEQ_OUT          (GT4_RXCHANBONDSEQ_OUT),
        .GT4_RXCHBONDEN_IN              (GT4_RXCHBONDEN_IN),
        .GT4_RXCHBONDLEVEL_IN           (GT4_RXCHBONDLEVEL_IN),
        .GT4_RXCHBONDMASTER_IN          (GT4_RXCHBONDMASTER_IN),
        .GT4_RXCHBONDO_OUT              (GT4_RXCHBONDO_OUT),
        .GT4_RXCHBONDSLAVE_IN           (GT4_RXCHBONDSLAVE_IN),
        //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
        .GT4_RXCHANISALIGNED_OUT        (GT4_RXCHANISALIGNED_OUT),
        .GT4_RXCHANREALIGN_OUT          (GT4_RXCHANREALIGN_OUT),
        //------------------ Receive Ports - RX Equailizer Ports -------------------
        .GT4_RXLPMHFHOLD_IN             (gt4_rxlpmhfhold_i),
        .GT4_RXLPMLFHOLD_IN             (gt4_rxlpmlfhold_i),
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .GT4_RXOUTCLK_OUT               (gt4_rxoutclk_i),
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .GT4_GTRXRESET_IN               (gt4_gtrxreset_i),
        .GT4_RXPMARESET_IN              (GT4_RXPMARESET_IN),
        //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        .GT4_RXCHARISK_OUT              (GT4_RXCHARISK_OUT),
        //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
        .GT4_RXCHBONDI_IN               (GT4_RXCHBONDI_IN),
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .GT4_RXRESETDONE_OUT            (gt4_rxresetdone_i),
        //------------------- TX Initialization and Reset Ports --------------------
        .GT4_GTTXRESET_IN               (gt4_gttxreset_i),
        .GT4_TXUSERRDY_IN               (gt4_txuserrdy_i),
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .GT4_TXUSRCLK_IN                (GT4_TXUSRCLK_IN),
        .GT4_TXUSRCLK2_IN               (GT4_TXUSRCLK2_IN),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .GT4_TXDATA_IN                  (GT4_TXDATA_IN),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .GT4_GTXTXN_OUT                 (GT4_GTXTXN_OUT),
        .GT4_GTXTXP_OUT                 (GT4_GTXTXP_OUT),
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .GT4_TXOUTCLK_OUT               (GT4_TXOUTCLK_OUT),
        .GT4_TXOUTCLKFABRIC_OUT         (GT4_TXOUTCLKFABRIC_OUT),
        .GT4_TXOUTCLKPCS_OUT            (GT4_TXOUTCLKPCS_OUT),
        //------------------- Transmit Ports - TX Gearbox Ports --------------------
        .GT4_TXCHARISK_IN               (GT4_TXCHARISK_IN),
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .GT4_TXRESETDONE_OUT            (gt4_txresetdone_i),


  
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT5  (X1Y9)

        //------------------------------- CPLL Ports -------------------------------
        .GT5_CPLLFBCLKLOST_OUT          (GT5_CPLLFBCLKLOST_OUT),
        .GT5_CPLLLOCK_OUT               (gt5_cplllock_i),
        .GT5_CPLLLOCKDETCLK_IN          (GT5_CPLLLOCKDETCLK_IN),
        .GT5_CPLLREFCLKLOST_OUT         (gt5_cpllrefclklost_i),
        .GT5_CPLLRESET_IN               (gt5_cpllreset_i),
        //------------------------ Channel - Clocking Ports ------------------------
        .GT5_GTREFCLK0_IN               (GT5_GTREFCLK0_IN),
        //-------------------------- Channel - DRP Ports  --------------------------
        .GT5_DRPADDR_IN                 (GT5_DRPADDR_IN),
        .GT5_DRPCLK_IN                  (GT5_DRPCLK_IN),
        .GT5_DRPDI_IN                   (GT5_DRPDI_IN),
        .GT5_DRPDO_OUT                  (GT5_DRPDO_OUT),
        .GT5_DRPEN_IN                   (GT5_DRPEN_IN),
        .GT5_DRPRDY_OUT                 (GT5_DRPRDY_OUT),
        .GT5_DRPWE_IN                   (GT5_DRPWE_IN),
        //----------------------------- Loopback Ports -----------------------------
        .GT5_LOOPBACK_IN                (GT5_LOOPBACK_IN),
        //------------------- RX Initialization and Reset Ports --------------------
        .GT5_RXUSERRDY_IN               (gt5_rxuserrdy_i),
        //------------------------ RX Margin Analysis Ports ------------------------
        .GT5_EYESCANDATAERROR_OUT       (GT5_EYESCANDATAERROR_OUT),
        //----------------------- Receive Ports - CDR Ports ------------------------
        .GT5_RXCDRLOCK_OUT              (GT5_RXCDRLOCK_OUT),
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .GT5_RXUSRCLK_IN                (GT5_RXUSRCLK_IN),
        .GT5_RXUSRCLK2_IN               (GT5_RXUSRCLK2_IN),
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .GT5_RXDATA_OUT                 (GT5_RXDATA_OUT),
        //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
        .GT5_RXDISPERR_OUT              (GT5_RXDISPERR_OUT),
        .GT5_RXNOTINTABLE_OUT           (GT5_RXNOTINTABLE_OUT),
        //------------------------- Receive Ports - RX AFE -------------------------
        .GT5_GTXRXP_IN                  (GT5_GTXRXP_IN),
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .GT5_GTXRXN_IN                  (GT5_GTXRXN_IN),
        //---------------- Receive Ports - RX Channel Bonding Ports ----------------
        .GT5_RXCHANBONDSEQ_OUT          (GT5_RXCHANBONDSEQ_OUT),
        .GT5_RXCHBONDEN_IN              (GT5_RXCHBONDEN_IN),
        .GT5_RXCHBONDLEVEL_IN           (GT5_RXCHBONDLEVEL_IN),
        .GT5_RXCHBONDMASTER_IN          (GT5_RXCHBONDMASTER_IN),
        .GT5_RXCHBONDO_OUT              (GT5_RXCHBONDO_OUT),
        .GT5_RXCHBONDSLAVE_IN           (GT5_RXCHBONDSLAVE_IN),
        //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
        .GT5_RXCHANISALIGNED_OUT        (GT5_RXCHANISALIGNED_OUT),
        .GT5_RXCHANREALIGN_OUT          (GT5_RXCHANREALIGN_OUT),
        //------------------ Receive Ports - RX Equailizer Ports -------------------
        .GT5_RXLPMHFHOLD_IN             (gt5_rxlpmhfhold_i),
        .GT5_RXLPMLFHOLD_IN             (gt5_rxlpmlfhold_i),
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .GT5_RXOUTCLK_OUT               (gt5_rxoutclk_i),
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .GT5_GTRXRESET_IN               (gt5_gtrxreset_i),
        .GT5_RXPMARESET_IN              (GT5_RXPMARESET_IN),
        //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        .GT5_RXCHARISK_OUT              (GT5_RXCHARISK_OUT),
        //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
        .GT5_RXCHBONDI_IN               (GT5_RXCHBONDI_IN),
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .GT5_RXRESETDONE_OUT            (gt5_rxresetdone_i),
        //------------------- TX Initialization and Reset Ports --------------------
        .GT5_GTTXRESET_IN               (gt5_gttxreset_i),
        .GT5_TXUSERRDY_IN               (gt5_txuserrdy_i),
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .GT5_TXUSRCLK_IN                (GT5_TXUSRCLK_IN),
        .GT5_TXUSRCLK2_IN               (GT5_TXUSRCLK2_IN),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .GT5_TXDATA_IN                  (GT5_TXDATA_IN),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .GT5_GTXTXN_OUT                 (GT5_GTXTXN_OUT),
        .GT5_GTXTXP_OUT                 (GT5_GTXTXP_OUT),
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .GT5_TXOUTCLK_OUT               (GT5_TXOUTCLK_OUT),
        .GT5_TXOUTCLKFABRIC_OUT         (GT5_TXOUTCLKFABRIC_OUT),
        .GT5_TXOUTCLKPCS_OUT            (GT5_TXOUTCLKPCS_OUT),
        //------------------- Transmit Ports - TX Gearbox Ports --------------------
        .GT5_TXCHARISK_IN               (GT5_TXCHARISK_IN),
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .GT5_TXRESETDONE_OUT            (gt5_txresetdone_i),


  
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT6  (X1Y10)

        //------------------------------- CPLL Ports -------------------------------
        .GT6_CPLLFBCLKLOST_OUT          (GT6_CPLLFBCLKLOST_OUT),
        .GT6_CPLLLOCK_OUT               (gt6_cplllock_i),
        .GT6_CPLLLOCKDETCLK_IN          (GT6_CPLLLOCKDETCLK_IN),
        .GT6_CPLLREFCLKLOST_OUT         (gt6_cpllrefclklost_i),
        .GT6_CPLLRESET_IN               (gt6_cpllreset_i),
        //------------------------ Channel - Clocking Ports ------------------------
        .GT6_GTREFCLK0_IN               (GT6_GTREFCLK0_IN),
        //-------------------------- Channel - DRP Ports  --------------------------
        .GT6_DRPADDR_IN                 (GT6_DRPADDR_IN),
        .GT6_DRPCLK_IN                  (GT6_DRPCLK_IN),
        .GT6_DRPDI_IN                   (GT6_DRPDI_IN),
        .GT6_DRPDO_OUT                  (GT6_DRPDO_OUT),
        .GT6_DRPEN_IN                   (GT6_DRPEN_IN),
        .GT6_DRPRDY_OUT                 (GT6_DRPRDY_OUT),
        .GT6_DRPWE_IN                   (GT6_DRPWE_IN),
        //----------------------------- Loopback Ports -----------------------------
        .GT6_LOOPBACK_IN                (GT6_LOOPBACK_IN),
        //------------------- RX Initialization and Reset Ports --------------------
        .GT6_RXUSERRDY_IN               (gt6_rxuserrdy_i),
        //------------------------ RX Margin Analysis Ports ------------------------
        .GT6_EYESCANDATAERROR_OUT       (GT6_EYESCANDATAERROR_OUT),
        //----------------------- Receive Ports - CDR Ports ------------------------
        .GT6_RXCDRLOCK_OUT              (GT6_RXCDRLOCK_OUT),
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .GT6_RXUSRCLK_IN                (GT6_RXUSRCLK_IN),
        .GT6_RXUSRCLK2_IN               (GT6_RXUSRCLK2_IN),
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .GT6_RXDATA_OUT                 (GT6_RXDATA_OUT),
        //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
        .GT6_RXDISPERR_OUT              (GT6_RXDISPERR_OUT),
        .GT6_RXNOTINTABLE_OUT           (GT6_RXNOTINTABLE_OUT),
        //------------------------- Receive Ports - RX AFE -------------------------
        .GT6_GTXRXP_IN                  (GT6_GTXRXP_IN),
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .GT6_GTXRXN_IN                  (GT6_GTXRXN_IN),
        //---------------- Receive Ports - RX Channel Bonding Ports ----------------
        .GT6_RXCHANBONDSEQ_OUT          (GT6_RXCHANBONDSEQ_OUT),
        .GT6_RXCHBONDEN_IN              (GT6_RXCHBONDEN_IN),
        .GT6_RXCHBONDLEVEL_IN           (GT6_RXCHBONDLEVEL_IN),
        .GT6_RXCHBONDMASTER_IN          (GT6_RXCHBONDMASTER_IN),
        .GT6_RXCHBONDO_OUT              (GT6_RXCHBONDO_OUT),
        .GT6_RXCHBONDSLAVE_IN           (GT6_RXCHBONDSLAVE_IN),
        //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
        .GT6_RXCHANISALIGNED_OUT        (GT6_RXCHANISALIGNED_OUT),
        .GT6_RXCHANREALIGN_OUT          (GT6_RXCHANREALIGN_OUT),
        //------------------ Receive Ports - RX Equailizer Ports -------------------
        .GT6_RXLPMHFHOLD_IN             (gt6_rxlpmhfhold_i),
        .GT6_RXLPMLFHOLD_IN             (gt6_rxlpmlfhold_i),
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .GT6_RXOUTCLK_OUT               (gt6_rxoutclk_i),
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .GT6_GTRXRESET_IN               (gt6_gtrxreset_i),
        .GT6_RXPMARESET_IN              (GT6_RXPMARESET_IN),
        //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        .GT6_RXCHARISK_OUT              (GT6_RXCHARISK_OUT),
        //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
        .GT6_RXCHBONDI_IN               (GT6_RXCHBONDI_IN),
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .GT6_RXRESETDONE_OUT            (gt6_rxresetdone_i),
        //------------------- TX Initialization and Reset Ports --------------------
        .GT6_GTTXRESET_IN               (gt6_gttxreset_i),
        .GT6_TXUSERRDY_IN               (gt6_txuserrdy_i),
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .GT6_TXUSRCLK_IN                (GT6_TXUSRCLK_IN),
        .GT6_TXUSRCLK2_IN               (GT6_TXUSRCLK2_IN),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .GT6_TXDATA_IN                  (GT6_TXDATA_IN),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .GT6_GTXTXN_OUT                 (GT6_GTXTXN_OUT),
        .GT6_GTXTXP_OUT                 (GT6_GTXTXP_OUT),
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .GT6_TXOUTCLK_OUT               (GT6_TXOUTCLK_OUT),
        .GT6_TXOUTCLKFABRIC_OUT         (GT6_TXOUTCLKFABRIC_OUT),
        .GT6_TXOUTCLKPCS_OUT            (GT6_TXOUTCLKPCS_OUT),
        //------------------- Transmit Ports - TX Gearbox Ports --------------------
        .GT6_TXCHARISK_IN               (GT6_TXCHARISK_IN),
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .GT6_TXRESETDONE_OUT            (gt6_txresetdone_i),


  
        //_____________________________________________________________________
        //_____________________________________________________________________
        //GT7  (X1Y11)

        //------------------------------- CPLL Ports -------------------------------
        .GT7_CPLLFBCLKLOST_OUT          (GT7_CPLLFBCLKLOST_OUT),
        .GT7_CPLLLOCK_OUT               (gt7_cplllock_i),
        .GT7_CPLLLOCKDETCLK_IN          (GT7_CPLLLOCKDETCLK_IN),
        .GT7_CPLLREFCLKLOST_OUT         (gt7_cpllrefclklost_i),
        .GT7_CPLLRESET_IN               (gt7_cpllreset_i),
        //------------------------ Channel - Clocking Ports ------------------------
        .GT7_GTREFCLK0_IN               (GT7_GTREFCLK0_IN),
        //-------------------------- Channel - DRP Ports  --------------------------
        .GT7_DRPADDR_IN                 (GT7_DRPADDR_IN),
        .GT7_DRPCLK_IN                  (GT7_DRPCLK_IN),
        .GT7_DRPDI_IN                   (GT7_DRPDI_IN),
        .GT7_DRPDO_OUT                  (GT7_DRPDO_OUT),
        .GT7_DRPEN_IN                   (GT7_DRPEN_IN),
        .GT7_DRPRDY_OUT                 (GT7_DRPRDY_OUT),
        .GT7_DRPWE_IN                   (GT7_DRPWE_IN),
        //----------------------------- Loopback Ports -----------------------------
        .GT7_LOOPBACK_IN                (GT7_LOOPBACK_IN),
        //------------------- RX Initialization and Reset Ports --------------------
        .GT7_RXUSERRDY_IN               (gt7_rxuserrdy_i),
        //------------------------ RX Margin Analysis Ports ------------------------
        .GT7_EYESCANDATAERROR_OUT       (GT7_EYESCANDATAERROR_OUT),
        //----------------------- Receive Ports - CDR Ports ------------------------
        .GT7_RXCDRLOCK_OUT              (GT7_RXCDRLOCK_OUT),
        //---------------- Receive Ports - FPGA RX Interface Ports -----------------
        .GT7_RXUSRCLK_IN                (GT7_RXUSRCLK_IN),
        .GT7_RXUSRCLK2_IN               (GT7_RXUSRCLK2_IN),
        //---------------- Receive Ports - FPGA RX interface Ports -----------------
        .GT7_RXDATA_OUT                 (GT7_RXDATA_OUT),
        //---------------- Receive Ports - RX 8B/10B Decoder Ports -----------------
        .GT7_RXDISPERR_OUT              (GT7_RXDISPERR_OUT),
        .GT7_RXNOTINTABLE_OUT           (GT7_RXNOTINTABLE_OUT),
        //------------------------- Receive Ports - RX AFE -------------------------
        .GT7_GTXRXP_IN                  (GT7_GTXRXP_IN),
        //---------------------- Receive Ports - RX AFE Ports ----------------------
        .GT7_GTXRXN_IN                  (GT7_GTXRXN_IN),
        //---------------- Receive Ports - RX Channel Bonding Ports ----------------
        .GT7_RXCHANBONDSEQ_OUT          (GT7_RXCHANBONDSEQ_OUT),
        .GT7_RXCHBONDEN_IN              (GT7_RXCHBONDEN_IN),
        .GT7_RXCHBONDLEVEL_IN           (GT7_RXCHBONDLEVEL_IN),
        .GT7_RXCHBONDMASTER_IN          (GT7_RXCHBONDMASTER_IN),
        .GT7_RXCHBONDO_OUT              (GT7_RXCHBONDO_OUT),
        .GT7_RXCHBONDSLAVE_IN           (GT7_RXCHBONDSLAVE_IN),
        //--------------- Receive Ports - RX Channel Bonding Ports  ----------------
        .GT7_RXCHANISALIGNED_OUT        (GT7_RXCHANISALIGNED_OUT),
        .GT7_RXCHANREALIGN_OUT          (GT7_RXCHANREALIGN_OUT),
        //------------------ Receive Ports - RX Equailizer Ports -------------------
        .GT7_RXLPMHFHOLD_IN             (gt7_rxlpmhfhold_i),
        .GT7_RXLPMLFHOLD_IN             (gt7_rxlpmlfhold_i),
        //------------- Receive Ports - RX Fabric Output Control Ports -------------
        .GT7_RXOUTCLK_OUT               (gt7_rxoutclk_i),
        //----------- Receive Ports - RX Initialization and Reset Ports ------------
        .GT7_GTRXRESET_IN               (gt7_gtrxreset_i),
        .GT7_RXPMARESET_IN              (GT7_RXPMARESET_IN),
        //----------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        .GT7_RXCHARISK_OUT              (GT7_RXCHARISK_OUT),
        //---------------- Receive Ports - Rx Channel Bonding Ports ----------------
        .GT7_RXCHBONDI_IN               (GT7_RXCHBONDI_IN),
        //------------ Receive Ports -RX Initialization and Reset Ports ------------
        .GT7_RXRESETDONE_OUT            (gt7_rxresetdone_i),
        //------------------- TX Initialization and Reset Ports --------------------
        .GT7_GTTXRESET_IN               (gt7_gttxreset_i),
        .GT7_TXUSERRDY_IN               (gt7_txuserrdy_i),
        //---------------- Transmit Ports - FPGA TX Interface Ports ----------------
        .GT7_TXUSRCLK_IN                (GT7_TXUSRCLK_IN),
        .GT7_TXUSRCLK2_IN               (GT7_TXUSRCLK2_IN),
        //---------------- Transmit Ports - TX Data Path interface -----------------
        .GT7_TXDATA_IN                  (GT7_TXDATA_IN),
        //-------------- Transmit Ports - TX Driver and OOB signaling --------------
        .GT7_GTXTXN_OUT                 (GT7_GTXTXN_OUT),
        .GT7_GTXTXP_OUT                 (GT7_GTXTXP_OUT),
        //--------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        .GT7_TXOUTCLK_OUT               (GT7_TXOUTCLK_OUT),
        .GT7_TXOUTCLKFABRIC_OUT         (GT7_TXOUTCLKFABRIC_OUT),
        .GT7_TXOUTCLKPCS_OUT            (GT7_TXOUTCLKPCS_OUT),
        //------------------- Transmit Ports - TX Gearbox Ports --------------------
        .GT7_TXCHARISK_IN               (GT7_TXCHARISK_IN),
        //----------- Transmit Ports - TX Initialization and Reset Ports -----------
        .GT7_TXRESETDONE_OUT            (gt7_txresetdone_i),




    //____________________________COMMON PORTS________________________________
        //-------------------- Common Block  - Ref Clock Ports ---------------------
        .GT0_GTREFCLK0_COMMON_IN        (GT0_GTREFCLK0_COMMON_IN),
        //----------------------- Common Block - QPLL Ports ------------------------
        .GT0_QPLLLOCK_OUT               (gt0_qplllock_i),
        .GT0_QPLLLOCKDETCLK_IN          (GT0_QPLLLOCKDETCLK_IN),
        .GT0_QPLLREFCLKLOST_OUT         (gt0_qpllrefclklost_i),
        .GT0_QPLLRESET_IN               (gt0_qpllreset_i),


    //____________________________COMMON PORTS________________________________
        //-------------------- Common Block  - Ref Clock Ports ---------------------
        .GT1_GTREFCLK0_COMMON_IN        (GT1_GTREFCLK0_COMMON_IN),
        //----------------------- Common Block - QPLL Ports ------------------------
        .GT1_QPLLLOCK_OUT               (gt1_qplllock_i),
        .GT1_QPLLLOCKDETCLK_IN          (GT1_QPLLLOCKDETCLK_IN),
        .GT1_QPLLREFCLKLOST_OUT         (gt1_qpllrefclklost_i),
        .GT1_QPLLRESET_IN               (gt1_qpllreset_i)

    );


    assign  gt0_rxdfelpmreset_i                  =  tied_to_ground_i;
    assign  gt1_rxdfelpmreset_i                  =  tied_to_ground_i;
    assign  gt2_rxdfelpmreset_i                  =  tied_to_ground_i;
    assign  gt3_rxdfelpmreset_i                  =  tied_to_ground_i;
    assign  gt4_rxdfelpmreset_i                  =  tied_to_ground_i;
    assign  gt5_rxdfelpmreset_i                  =  tied_to_ground_i;
    assign  gt6_rxdfelpmreset_i                  =  tied_to_ground_i;
    assign  gt7_rxdfelpmreset_i                  =  tied_to_ground_i;


    assign  GT0_CPLLLOCK_OUT                     =  gt0_cplllock_i;
    assign  GT0_TXRESETDONE_OUT                  =  gt0_txresetdone_i;
    assign  GT0_RXRESETDONE_OUT                  =  gt0_rxresetdone_i;
    assign  GT1_CPLLLOCK_OUT                     =  gt1_cplllock_i;
    assign  GT1_TXRESETDONE_OUT                  =  gt1_txresetdone_i;
    assign  GT1_RXRESETDONE_OUT                  =  gt1_rxresetdone_i;
    assign  GT2_CPLLLOCK_OUT                     =  gt2_cplllock_i;
    assign  GT2_TXRESETDONE_OUT                  =  gt2_txresetdone_i;
    assign  GT2_RXRESETDONE_OUT                  =  gt2_rxresetdone_i;
    assign  GT3_CPLLLOCK_OUT                     =  gt3_cplllock_i;
    assign  GT3_TXRESETDONE_OUT                  =  gt3_txresetdone_i;
    assign  GT3_RXRESETDONE_OUT                  =  gt3_rxresetdone_i;
    assign  GT4_CPLLLOCK_OUT                     =  gt4_cplllock_i;
    assign  GT4_TXRESETDONE_OUT                  =  gt4_txresetdone_i;
    assign  GT4_RXRESETDONE_OUT                  =  gt4_rxresetdone_i;
    assign  GT5_CPLLLOCK_OUT                     =  gt5_cplllock_i;
    assign  GT5_TXRESETDONE_OUT                  =  gt5_txresetdone_i;
    assign  GT5_RXRESETDONE_OUT                  =  gt5_rxresetdone_i;
    assign  GT6_CPLLLOCK_OUT                     =  gt6_cplllock_i;
    assign  GT6_TXRESETDONE_OUT                  =  gt6_txresetdone_i;
    assign  GT6_RXRESETDONE_OUT                  =  gt6_rxresetdone_i;
    assign  GT7_CPLLLOCK_OUT                     =  gt7_cplllock_i;
    assign  GT7_TXRESETDONE_OUT                  =  gt7_txresetdone_i;
    assign  GT7_RXRESETDONE_OUT                  =  gt7_rxresetdone_i;
    assign  GT0_QPLLLOCK_OUT                     =  gt0_qplllock_i;
    assign  GT1_QPLLLOCK_OUT                     =  gt1_qplllock_i;

generate
if (EXAMPLE_USE_CHIPSCOPE == 1) 
begin : chipscope
    assign  gt0_cpllreset_i                      =  GT0_CPLLRESET_IN || gt0_cpllreset_t;
    assign  gt0_gttxreset_i                      =  GT0_GTTXRESET_IN || gt0_gttxreset_t;
    assign  gt0_gtrxreset_i                      =  GT0_GTRXRESET_IN || gt0_gtrxreset_t;
    assign  gt0_txuserrdy_i                      =  GT0_TXUSERRDY_IN || gt0_txuserrdy_t;
    assign  gt0_rxuserrdy_i                      =  GT0_RXUSERRDY_IN || gt0_rxuserrdy_t;
    assign  gt1_cpllreset_i                      =  GT1_CPLLRESET_IN || gt1_cpllreset_t;
    assign  gt1_gttxreset_i                      =  GT1_GTTXRESET_IN || gt1_gttxreset_t;
    assign  gt1_gtrxreset_i                      =  GT1_GTRXRESET_IN || gt1_gtrxreset_t;
    assign  gt1_txuserrdy_i                      =  GT1_TXUSERRDY_IN || gt1_txuserrdy_t;
    assign  gt1_rxuserrdy_i                      =  GT1_RXUSERRDY_IN || gt1_rxuserrdy_t;
    assign  gt2_cpllreset_i                      =  GT2_CPLLRESET_IN || gt2_cpllreset_t;
    assign  gt2_gttxreset_i                      =  GT2_GTTXRESET_IN || gt2_gttxreset_t;
    assign  gt2_gtrxreset_i                      =  GT2_GTRXRESET_IN || gt2_gtrxreset_t;
    assign  gt2_txuserrdy_i                      =  GT2_TXUSERRDY_IN || gt2_txuserrdy_t;
    assign  gt2_rxuserrdy_i                      =  GT2_RXUSERRDY_IN || gt2_rxuserrdy_t;
    assign  gt3_cpllreset_i                      =  GT3_CPLLRESET_IN || gt3_cpllreset_t;
    assign  gt3_gttxreset_i                      =  GT3_GTTXRESET_IN || gt3_gttxreset_t;
    assign  gt3_gtrxreset_i                      =  GT3_GTRXRESET_IN || gt3_gtrxreset_t;
    assign  gt3_txuserrdy_i                      =  GT3_TXUSERRDY_IN || gt3_txuserrdy_t;
    assign  gt3_rxuserrdy_i                      =  GT3_RXUSERRDY_IN || gt3_rxuserrdy_t;
    assign  gt4_cpllreset_i                      =  GT4_CPLLRESET_IN || gt4_cpllreset_t;
    assign  gt4_gttxreset_i                      =  GT4_GTTXRESET_IN || gt4_gttxreset_t;
    assign  gt4_gtrxreset_i                      =  GT4_GTRXRESET_IN || gt4_gtrxreset_t;
    assign  gt4_txuserrdy_i                      =  GT4_TXUSERRDY_IN || gt4_txuserrdy_t;
    assign  gt4_rxuserrdy_i                      =  GT4_RXUSERRDY_IN || gt4_rxuserrdy_t;
    assign  gt5_cpllreset_i                      =  GT5_CPLLRESET_IN || gt5_cpllreset_t;
    assign  gt5_gttxreset_i                      =  GT5_GTTXRESET_IN || gt5_gttxreset_t;
    assign  gt5_gtrxreset_i                      =  GT5_GTRXRESET_IN || gt5_gtrxreset_t;
    assign  gt5_txuserrdy_i                      =  GT5_TXUSERRDY_IN || gt5_txuserrdy_t;
    assign  gt5_rxuserrdy_i                      =  GT5_RXUSERRDY_IN || gt5_rxuserrdy_t;
    assign  gt6_cpllreset_i                      =  GT6_CPLLRESET_IN || gt6_cpllreset_t;
    assign  gt6_gttxreset_i                      =  GT6_GTTXRESET_IN || gt6_gttxreset_t;
    assign  gt6_gtrxreset_i                      =  GT6_GTRXRESET_IN || gt6_gtrxreset_t;
    assign  gt6_txuserrdy_i                      =  GT6_TXUSERRDY_IN || gt6_txuserrdy_t;
    assign  gt6_rxuserrdy_i                      =  GT6_RXUSERRDY_IN || gt6_rxuserrdy_t;
    assign  gt7_cpllreset_i                      =  GT7_CPLLRESET_IN || gt7_cpllreset_t;
    assign  gt7_gttxreset_i                      =  GT7_GTTXRESET_IN || gt7_gttxreset_t;
    assign  gt7_gtrxreset_i                      =  GT7_GTRXRESET_IN || gt7_gtrxreset_t;
    assign  gt7_txuserrdy_i                      =  GT7_TXUSERRDY_IN || gt7_txuserrdy_t;
    assign  gt7_rxuserrdy_i                      =  GT7_RXUSERRDY_IN || gt7_rxuserrdy_t;
    assign  gt0_qpllreset_i                      =  GT0_QPLLRESET_IN || gt0_qpllreset_t;
    assign  gt1_qpllreset_i                      =  GT1_QPLLRESET_IN || gt1_qpllreset_t;
end
endgenerate 

generate
if (EXAMPLE_USE_CHIPSCOPE == 0) 
begin : no_chipscope
    assign  gt0_cpllreset_i                      =  gt0_cpllreset_t;
    assign  gt0_gttxreset_i                      =  gt0_gttxreset_t;
    assign  gt0_gtrxreset_i                      =  gt0_gtrxreset_t;
    assign  gt0_txuserrdy_i                      =  gt0_txuserrdy_t;
    assign  gt0_rxuserrdy_i                      =  gt0_rxuserrdy_t;
    assign  gt1_cpllreset_i                      =  gt1_cpllreset_t;
    assign  gt1_gttxreset_i                      =  gt1_gttxreset_t;
    assign  gt1_gtrxreset_i                      =  gt1_gtrxreset_t;
    assign  gt1_txuserrdy_i                      =  gt1_txuserrdy_t;
    assign  gt1_rxuserrdy_i                      =  gt1_rxuserrdy_t;
    assign  gt2_cpllreset_i                      =  gt2_cpllreset_t;
    assign  gt2_gttxreset_i                      =  gt2_gttxreset_t;
    assign  gt2_gtrxreset_i                      =  gt2_gtrxreset_t;
    assign  gt2_txuserrdy_i                      =  gt2_txuserrdy_t;
    assign  gt2_rxuserrdy_i                      =  gt2_rxuserrdy_t;
    assign  gt3_cpllreset_i                      =  gt3_cpllreset_t;
    assign  gt3_gttxreset_i                      =  gt3_gttxreset_t;
    assign  gt3_gtrxreset_i                      =  gt3_gtrxreset_t;
    assign  gt3_txuserrdy_i                      =  gt3_txuserrdy_t;
    assign  gt3_rxuserrdy_i                      =  gt3_rxuserrdy_t;
    assign  gt4_cpllreset_i                      =  gt4_cpllreset_t;
    assign  gt4_gttxreset_i                      =  gt4_gttxreset_t;
    assign  gt4_gtrxreset_i                      =  gt4_gtrxreset_t;
    assign  gt4_txuserrdy_i                      =  gt4_txuserrdy_t;
    assign  gt4_rxuserrdy_i                      =  gt4_rxuserrdy_t;
    assign  gt5_cpllreset_i                      =  gt5_cpllreset_t;
    assign  gt5_gttxreset_i                      =  gt5_gttxreset_t;
    assign  gt5_gtrxreset_i                      =  gt5_gtrxreset_t;
    assign  gt5_txuserrdy_i                      =  gt5_txuserrdy_t;
    assign  gt5_rxuserrdy_i                      =  gt5_rxuserrdy_t;
    assign  gt6_cpllreset_i                      =  gt6_cpllreset_t;
    assign  gt6_gttxreset_i                      =  gt6_gttxreset_t;
    assign  gt6_gtrxreset_i                      =  gt6_gtrxreset_t;
    assign  gt6_txuserrdy_i                      =  gt6_txuserrdy_t;
    assign  gt6_rxuserrdy_i                      =  gt6_rxuserrdy_t;
    assign  gt7_cpllreset_i                      =  gt7_cpllreset_t;
    assign  gt7_gttxreset_i                      =  gt7_gttxreset_t;
    assign  gt7_gtrxreset_i                      =  gt7_gtrxreset_t;
    assign  gt7_txuserrdy_i                      =  gt7_txuserrdy_t;
    assign  gt7_rxuserrdy_i                      =  gt7_rxuserrdy_t;
    assign  gt0_qpllreset_i                      =  gt0_qpllreset_t;
    assign  gt1_qpllreset_i                      =  gt1_qpllreset_t;
end
endgenerate 


serdes_coe_TX_STARTUP_FSM #
          (
           .GT_TYPE                  ("GTX"), //GTX or GTH or GTP
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("FALSE"),                       // the TX and RX Reset FSMs must
           .RX_QPLL_USED             ("FALSE"),                       // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt0_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (SYSCLK_IN),
        .TXUSERCLK                      (GT0_TXUSRCLK_IN),
        .SOFT_RESET                     (SOFT_RESET_IN),
        .QPLLREFCLKLOST                 (tied_to_ground_i),
        .CPLLREFCLKLOST                 (gt0_cpllrefclklost_i),
        .QPLLLOCK                       (tied_to_vcc_i),
        .CPLLLOCK                       (gt0_cplllock_i),
        .TXRESETDONE                    (gt0_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt0_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (gt0_cpllreset_t),
        .TX_FSM_RESET_DONE              (GT0_TX_FSM_RESET_DONE_OUT),
        .TXUSERRDY                      (gt0_txuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RETRY_COUNTER                  ()
           );


serdes_coe_TX_STARTUP_FSM #
          (
           .GT_TYPE                  ("GTX"), //GTX or GTH or GTP
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("FALSE"),                       // the TX and RX Reset FSMs must
           .RX_QPLL_USED             ("FALSE"),                       // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt1_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (SYSCLK_IN),
        .TXUSERCLK                      (GT1_TXUSRCLK_IN),
        .SOFT_RESET                     (SOFT_RESET_IN),
        .QPLLREFCLKLOST                 (tied_to_ground_i),
        .CPLLREFCLKLOST                 (gt1_cpllrefclklost_i),
        .QPLLLOCK                       (tied_to_vcc_i),
        .CPLLLOCK                       (gt1_cplllock_i),
        .TXRESETDONE                    (gt1_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt1_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (gt1_cpllreset_t),
        .TX_FSM_RESET_DONE              (GT1_TX_FSM_RESET_DONE_OUT),
        .TXUSERRDY                      (gt1_txuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RETRY_COUNTER                  ()
           );


serdes_coe_TX_STARTUP_FSM #
          (
           .GT_TYPE                  ("GTX"), //GTX or GTH or GTP
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("FALSE"),                       // the TX and RX Reset FSMs must
           .RX_QPLL_USED             ("FALSE"),                       // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt2_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (SYSCLK_IN),
        .TXUSERCLK                      (GT2_TXUSRCLK_IN),
        .SOFT_RESET                     (SOFT_RESET_IN),
        .QPLLREFCLKLOST                 (tied_to_ground_i),
        .CPLLREFCLKLOST                 (gt2_cpllrefclklost_i),
        .QPLLLOCK                       (tied_to_vcc_i),
        .CPLLLOCK                       (gt2_cplllock_i),
        .TXRESETDONE                    (gt2_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt2_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (gt2_cpllreset_t),
        .TX_FSM_RESET_DONE              (GT2_TX_FSM_RESET_DONE_OUT),
        .TXUSERRDY                      (gt2_txuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RETRY_COUNTER                  ()
           );


serdes_coe_TX_STARTUP_FSM #
          (
           .GT_TYPE                  ("GTX"), //GTX or GTH or GTP
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("FALSE"),                       // the TX and RX Reset FSMs must
           .RX_QPLL_USED             ("FALSE"),                       // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt3_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (SYSCLK_IN),
        .TXUSERCLK                      (GT3_TXUSRCLK_IN),
        .SOFT_RESET                     (SOFT_RESET_IN),
        .QPLLREFCLKLOST                 (tied_to_ground_i),
        .CPLLREFCLKLOST                 (gt3_cpllrefclklost_i),
        .QPLLLOCK                       (tied_to_vcc_i),
        .CPLLLOCK                       (gt3_cplllock_i),
        .TXRESETDONE                    (gt3_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt3_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (gt3_cpllreset_t),
        .TX_FSM_RESET_DONE              (GT3_TX_FSM_RESET_DONE_OUT),
        .TXUSERRDY                      (gt3_txuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RETRY_COUNTER                  ()
           );


serdes_coe_TX_STARTUP_FSM #
          (
           .GT_TYPE                  ("GTX"), //GTX or GTH or GTP
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("FALSE"),                       // the TX and RX Reset FSMs must
           .RX_QPLL_USED             ("FALSE"),                       // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt4_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (SYSCLK_IN),
        .TXUSERCLK                      (GT4_TXUSRCLK_IN),
        .SOFT_RESET                     (SOFT_RESET_IN),
        .QPLLREFCLKLOST                 (tied_to_ground_i),
        .CPLLREFCLKLOST                 (gt4_cpllrefclklost_i),
        .QPLLLOCK                       (tied_to_vcc_i),
        .CPLLLOCK                       (gt4_cplllock_i),
        .TXRESETDONE                    (gt4_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt4_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (gt4_cpllreset_t),
        .TX_FSM_RESET_DONE              (GT4_TX_FSM_RESET_DONE_OUT),
        .TXUSERRDY                      (gt4_txuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RETRY_COUNTER                  ()
           );


serdes_coe_TX_STARTUP_FSM #
          (
           .GT_TYPE                  ("GTX"), //GTX or GTH or GTP
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("FALSE"),                       // the TX and RX Reset FSMs must
           .RX_QPLL_USED             ("FALSE"),                       // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt5_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (SYSCLK_IN),
        .TXUSERCLK                      (GT5_TXUSRCLK_IN),
        .SOFT_RESET                     (SOFT_RESET_IN),
        .QPLLREFCLKLOST                 (tied_to_ground_i),
        .CPLLREFCLKLOST                 (gt5_cpllrefclklost_i),
        .QPLLLOCK                       (tied_to_vcc_i),
        .CPLLLOCK                       (gt5_cplllock_i),
        .TXRESETDONE                    (gt5_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt5_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (gt5_cpllreset_t),
        .TX_FSM_RESET_DONE              (GT5_TX_FSM_RESET_DONE_OUT),
        .TXUSERRDY                      (gt5_txuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RETRY_COUNTER                  ()
           );


serdes_coe_TX_STARTUP_FSM #
          (
           .GT_TYPE                  ("GTX"), //GTX or GTH or GTP
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("FALSE"),                       // the TX and RX Reset FSMs must
           .RX_QPLL_USED             ("FALSE"),                       // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt6_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (SYSCLK_IN),
        .TXUSERCLK                      (GT6_TXUSRCLK_IN),
        .SOFT_RESET                     (SOFT_RESET_IN),
        .QPLLREFCLKLOST                 (tied_to_ground_i),
        .CPLLREFCLKLOST                 (gt6_cpllrefclklost_i),
        .QPLLLOCK                       (tied_to_vcc_i),
        .CPLLLOCK                       (gt6_cplllock_i),
        .TXRESETDONE                    (gt6_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt6_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (gt6_cpllreset_t),
        .TX_FSM_RESET_DONE              (GT6_TX_FSM_RESET_DONE_OUT),
        .TXUSERRDY                      (gt6_txuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RETRY_COUNTER                  ()
           );


serdes_coe_TX_STARTUP_FSM #
          (
           .GT_TYPE                  ("GTX"), //GTX or GTH or GTP
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),           // Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("FALSE"),                       // the TX and RX Reset FSMs must
           .RX_QPLL_USED             ("FALSE"),                       // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")               // Decision if a manual phase-alignment is necessary or the automatic 
                                                                     // is enough. For single-lane applications the automatic alignment is 
                                                                     // sufficient              
             ) 
gt7_txresetfsm_i      
            ( 
        .STABLE_CLOCK                   (SYSCLK_IN),
        .TXUSERCLK                      (GT7_TXUSRCLK_IN),
        .SOFT_RESET                     (SOFT_RESET_IN),
        .QPLLREFCLKLOST                 (tied_to_ground_i),
        .CPLLREFCLKLOST                 (gt7_cpllrefclklost_i),
        .QPLLLOCK                       (tied_to_vcc_i),
        .CPLLLOCK                       (gt7_cplllock_i),
        .TXRESETDONE                    (gt7_txresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .GTTXRESET                      (gt7_gttxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (gt7_cpllreset_t),
        .TX_FSM_RESET_DONE              (GT7_TX_FSM_RESET_DONE_OUT),
        .TXUSERRDY                      (gt7_txuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RETRY_COUNTER                  ()
           );



serdes_coe_RX_STARTUP_FSM  #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .GT_TYPE                  ("GTX"), //GTX or GTH or GTP
           .EQ_MODE                  ("LPM"),                   //Rx Equalization Mode - Set to DFE or LPM
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),              //Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("FALSE"),                          // the TX and RX Reset FSMs must
           .RX_QPLL_USED             ("FALSE"),                          // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")                 // Decision if a manual phase-alignment is necessary or the automatic 
                                                                         // is enough. For single-lane applications the automatic alignment is 
                                                                         // sufficient              
             )     
gt0_rxresetfsm_i
             ( 
        .STABLE_CLOCK                   (SYSCLK_IN),
        .RXUSERCLK                      (GT0_RXUSRCLK_IN),
        .SOFT_RESET                     (SOFT_RESET_IN),
        .DONT_RESET_ON_DATA_ERROR       (DONT_RESET_ON_DATA_ERROR_IN),
        .QPLLREFCLKLOST                 (tied_to_ground_i),
        .CPLLREFCLKLOST                 (gt0_cpllrefclklost_i),
        .QPLLLOCK                       (tied_to_vcc_i),
        .CPLLLOCK                       (gt0_cplllock_i),
        .RXRESETDONE                    (gt0_rxresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .RECCLK_STABLE                  (gt0_recclk_stable_i),
        .RECCLK_MONITOR_RESTART         (tied_to_ground_i),
        .DATA_VALID                     (GT0_DATA_VALID_IN),
        .TXUSERRDY                      (gt0_txuserrdy_i),
        .GTRXRESET                      (gt0_gtrxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .RX_FSM_RESET_DONE              (GT0_RX_FSM_RESET_DONE_OUT),
        .RXUSERRDY                      (gt0_rxuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RXDFEAGCHOLD                   (gt0_rxdfeagchold_i),
        .RXDFELFHOLD                    (gt0_rxdfelfhold_i),
        .RXLPMLFHOLD                    (gt0_rxlpmlfhold_i),
        .RXLPMHFHOLD                    (gt0_rxlpmhfhold_i),
        .RETRY_COUNTER                  ()
           );

serdes_coe_RX_STARTUP_FSM  #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .GT_TYPE                  ("GTX"), //GTX or GTH or GTP
           .EQ_MODE                  ("LPM"),                   //Rx Equalization Mode - Set to DFE or LPM
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),              //Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("FALSE"),                          // the TX and RX Reset FSMs must
           .RX_QPLL_USED             ("FALSE"),                          // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")                 // Decision if a manual phase-alignment is necessary or the automatic 
                                                                         // is enough. For single-lane applications the automatic alignment is 
                                                                         // sufficient              
             )     
gt1_rxresetfsm_i
             ( 
        .STABLE_CLOCK                   (SYSCLK_IN),
        .RXUSERCLK                      (GT1_RXUSRCLK_IN),
        .SOFT_RESET                     (SOFT_RESET_IN),
        .DONT_RESET_ON_DATA_ERROR       (DONT_RESET_ON_DATA_ERROR_IN),
        .QPLLREFCLKLOST                 (tied_to_ground_i),
        .CPLLREFCLKLOST                 (gt1_cpllrefclklost_i),
        .QPLLLOCK                       (tied_to_vcc_i),
        .CPLLLOCK                       (gt1_cplllock_i),
        .RXRESETDONE                    (gt1_rxresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .RECCLK_STABLE                  (gt1_recclk_stable_i),
        .RECCLK_MONITOR_RESTART         (tied_to_ground_i),
        .DATA_VALID                     (GT1_DATA_VALID_IN),
        .TXUSERRDY                      (gt1_txuserrdy_i),
        .GTRXRESET                      (gt1_gtrxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .RX_FSM_RESET_DONE              (GT1_RX_FSM_RESET_DONE_OUT),
        .RXUSERRDY                      (gt1_rxuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RXDFEAGCHOLD                   (gt1_rxdfeagchold_i),
        .RXDFELFHOLD                    (gt1_rxdfelfhold_i),
        .RXLPMLFHOLD                    (gt1_rxlpmlfhold_i),
        .RXLPMHFHOLD                    (gt1_rxlpmhfhold_i),
        .RETRY_COUNTER                  ()
           );

serdes_coe_RX_STARTUP_FSM  #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .GT_TYPE                  ("GTX"), //GTX or GTH or GTP
           .EQ_MODE                  ("LPM"),                   //Rx Equalization Mode - Set to DFE or LPM
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),              //Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("FALSE"),                          // the TX and RX Reset FSMs must
           .RX_QPLL_USED             ("FALSE"),                          // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")                 // Decision if a manual phase-alignment is necessary or the automatic 
                                                                         // is enough. For single-lane applications the automatic alignment is 
                                                                         // sufficient              
             )     
gt2_rxresetfsm_i
             ( 
        .STABLE_CLOCK                   (SYSCLK_IN),
        .RXUSERCLK                      (GT2_RXUSRCLK_IN),
        .SOFT_RESET                     (SOFT_RESET_IN),
        .DONT_RESET_ON_DATA_ERROR       (DONT_RESET_ON_DATA_ERROR_IN),
        .QPLLREFCLKLOST                 (tied_to_ground_i),
        .CPLLREFCLKLOST                 (gt2_cpllrefclklost_i),
        .QPLLLOCK                       (tied_to_vcc_i),
        .CPLLLOCK                       (gt2_cplllock_i),
        .RXRESETDONE                    (gt2_rxresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .RECCLK_STABLE                  (gt2_recclk_stable_i),
        .RECCLK_MONITOR_RESTART         (tied_to_ground_i),
        .DATA_VALID                     (GT2_DATA_VALID_IN),
        .TXUSERRDY                      (gt2_txuserrdy_i),
        .GTRXRESET                      (gt2_gtrxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .RX_FSM_RESET_DONE              (GT2_RX_FSM_RESET_DONE_OUT),
        .RXUSERRDY                      (gt2_rxuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RXDFEAGCHOLD                   (gt2_rxdfeagchold_i),
        .RXDFELFHOLD                    (gt2_rxdfelfhold_i),
        .RXLPMLFHOLD                    (gt2_rxlpmlfhold_i),
        .RXLPMHFHOLD                    (gt2_rxlpmhfhold_i),
        .RETRY_COUNTER                  ()
           );

serdes_coe_RX_STARTUP_FSM  #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .GT_TYPE                  ("GTX"), //GTX or GTH or GTP
           .EQ_MODE                  ("LPM"),                   //Rx Equalization Mode - Set to DFE or LPM
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),              //Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("FALSE"),                          // the TX and RX Reset FSMs must
           .RX_QPLL_USED             ("FALSE"),                          // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")                 // Decision if a manual phase-alignment is necessary or the automatic 
                                                                         // is enough. For single-lane applications the automatic alignment is 
                                                                         // sufficient              
             )     
gt3_rxresetfsm_i
             ( 
        .STABLE_CLOCK                   (SYSCLK_IN),
        .RXUSERCLK                      (GT3_RXUSRCLK_IN),
        .SOFT_RESET                     (SOFT_RESET_IN),
        .DONT_RESET_ON_DATA_ERROR       (DONT_RESET_ON_DATA_ERROR_IN),
        .QPLLREFCLKLOST                 (tied_to_ground_i),
        .CPLLREFCLKLOST                 (gt3_cpllrefclklost_i),
        .QPLLLOCK                       (tied_to_vcc_i),
        .CPLLLOCK                       (gt3_cplllock_i),
        .RXRESETDONE                    (gt3_rxresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .RECCLK_STABLE                  (gt3_recclk_stable_i),
        .RECCLK_MONITOR_RESTART         (tied_to_ground_i),
        .DATA_VALID                     (GT3_DATA_VALID_IN),
        .TXUSERRDY                      (gt3_txuserrdy_i),
        .GTRXRESET                      (gt3_gtrxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .RX_FSM_RESET_DONE              (GT3_RX_FSM_RESET_DONE_OUT),
        .RXUSERRDY                      (gt3_rxuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RXDFEAGCHOLD                   (gt3_rxdfeagchold_i),
        .RXDFELFHOLD                    (gt3_rxdfelfhold_i),
        .RXLPMLFHOLD                    (gt3_rxlpmlfhold_i),
        .RXLPMHFHOLD                    (gt3_rxlpmhfhold_i),
        .RETRY_COUNTER                  ()
           );

serdes_coe_RX_STARTUP_FSM  #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .GT_TYPE                  ("GTX"), //GTX or GTH or GTP
           .EQ_MODE                  ("LPM"),                   //Rx Equalization Mode - Set to DFE or LPM
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),              //Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("FALSE"),                          // the TX and RX Reset FSMs must
           .RX_QPLL_USED             ("FALSE"),                          // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")                 // Decision if a manual phase-alignment is necessary or the automatic 
                                                                         // is enough. For single-lane applications the automatic alignment is 
                                                                         // sufficient              
             )     
gt4_rxresetfsm_i
             ( 
        .STABLE_CLOCK                   (SYSCLK_IN),
        .RXUSERCLK                      (GT4_RXUSRCLK_IN),
        .SOFT_RESET                     (SOFT_RESET_IN),
        .DONT_RESET_ON_DATA_ERROR       (DONT_RESET_ON_DATA_ERROR_IN),
        .QPLLREFCLKLOST                 (tied_to_ground_i),
        .CPLLREFCLKLOST                 (gt4_cpllrefclklost_i),
        .QPLLLOCK                       (tied_to_vcc_i),
        .CPLLLOCK                       (gt4_cplllock_i),
        .RXRESETDONE                    (gt4_rxresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .RECCLK_STABLE                  (gt4_recclk_stable_i),
        .RECCLK_MONITOR_RESTART         (tied_to_ground_i),
        .DATA_VALID                     (GT4_DATA_VALID_IN),
        .TXUSERRDY                      (gt4_txuserrdy_i),
        .GTRXRESET                      (gt4_gtrxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .RX_FSM_RESET_DONE              (GT4_RX_FSM_RESET_DONE_OUT),
        .RXUSERRDY                      (gt4_rxuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RXDFEAGCHOLD                   (gt4_rxdfeagchold_i),
        .RXDFELFHOLD                    (gt4_rxdfelfhold_i),
        .RXLPMLFHOLD                    (gt4_rxlpmlfhold_i),
        .RXLPMHFHOLD                    (gt4_rxlpmhfhold_i),
        .RETRY_COUNTER                  ()
           );

serdes_coe_RX_STARTUP_FSM  #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .GT_TYPE                  ("GTX"), //GTX or GTH or GTP
           .EQ_MODE                  ("LPM"),                   //Rx Equalization Mode - Set to DFE or LPM
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),              //Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("FALSE"),                          // the TX and RX Reset FSMs must
           .RX_QPLL_USED             ("FALSE"),                          // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")                 // Decision if a manual phase-alignment is necessary or the automatic 
                                                                         // is enough. For single-lane applications the automatic alignment is 
                                                                         // sufficient              
             )     
gt5_rxresetfsm_i
             ( 
        .STABLE_CLOCK                   (SYSCLK_IN),
        .RXUSERCLK                      (GT5_RXUSRCLK_IN),
        .SOFT_RESET                     (SOFT_RESET_IN),
        .DONT_RESET_ON_DATA_ERROR       (DONT_RESET_ON_DATA_ERROR_IN),
        .QPLLREFCLKLOST                 (tied_to_ground_i),
        .CPLLREFCLKLOST                 (gt5_cpllrefclklost_i),
        .QPLLLOCK                       (tied_to_vcc_i),
        .CPLLLOCK                       (gt5_cplllock_i),
        .RXRESETDONE                    (gt5_rxresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .RECCLK_STABLE                  (gt5_recclk_stable_i),
        .RECCLK_MONITOR_RESTART         (tied_to_ground_i),
        .DATA_VALID                     (GT5_DATA_VALID_IN),
        .TXUSERRDY                      (gt5_txuserrdy_i),
        .GTRXRESET                      (gt5_gtrxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .RX_FSM_RESET_DONE              (GT5_RX_FSM_RESET_DONE_OUT),
        .RXUSERRDY                      (gt5_rxuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RXDFEAGCHOLD                   (gt5_rxdfeagchold_i),
        .RXDFELFHOLD                    (gt5_rxdfelfhold_i),
        .RXLPMLFHOLD                    (gt5_rxlpmlfhold_i),
        .RXLPMHFHOLD                    (gt5_rxlpmhfhold_i),
        .RETRY_COUNTER                  ()
           );

serdes_coe_RX_STARTUP_FSM  #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .GT_TYPE                  ("GTX"), //GTX or GTH or GTP
           .EQ_MODE                  ("LPM"),                   //Rx Equalization Mode - Set to DFE or LPM
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),              //Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("FALSE"),                          // the TX and RX Reset FSMs must
           .RX_QPLL_USED             ("FALSE"),                          // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")                 // Decision if a manual phase-alignment is necessary or the automatic 
                                                                         // is enough. For single-lane applications the automatic alignment is 
                                                                         // sufficient              
             )     
gt6_rxresetfsm_i
             ( 
        .STABLE_CLOCK                   (SYSCLK_IN),
        .RXUSERCLK                      (GT6_RXUSRCLK_IN),
        .SOFT_RESET                     (SOFT_RESET_IN),
        .DONT_RESET_ON_DATA_ERROR       (DONT_RESET_ON_DATA_ERROR_IN),
        .QPLLREFCLKLOST                 (tied_to_ground_i),
        .CPLLREFCLKLOST                 (gt6_cpllrefclklost_i),
        .QPLLLOCK                       (tied_to_vcc_i),
        .CPLLLOCK                       (gt6_cplllock_i),
        .RXRESETDONE                    (gt6_rxresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .RECCLK_STABLE                  (gt6_recclk_stable_i),
        .RECCLK_MONITOR_RESTART         (tied_to_ground_i),
        .DATA_VALID                     (GT6_DATA_VALID_IN),
        .TXUSERRDY                      (gt6_txuserrdy_i),
        .GTRXRESET                      (gt6_gtrxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .RX_FSM_RESET_DONE              (GT6_RX_FSM_RESET_DONE_OUT),
        .RXUSERRDY                      (gt6_rxuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RXDFEAGCHOLD                   (gt6_rxdfeagchold_i),
        .RXDFELFHOLD                    (gt6_rxdfelfhold_i),
        .RXLPMLFHOLD                    (gt6_rxlpmlfhold_i),
        .RXLPMHFHOLD                    (gt6_rxlpmhfhold_i),
        .RETRY_COUNTER                  ()
           );

serdes_coe_RX_STARTUP_FSM  #
          (
           .EXAMPLE_SIMULATION       (EXAMPLE_SIMULATION),
           .GT_TYPE                  ("GTX"), //GTX or GTH or GTP
           .EQ_MODE                  ("LPM"),                   //Rx Equalization Mode - Set to DFE or LPM
           .STABLE_CLOCK_PERIOD      (STABLE_CLOCK_PERIOD),              //Period of the stable clock driving this state-machine, unit is [ns]
           .RETRY_COUNTER_BITWIDTH   (8), 
           .TX_QPLL_USED             ("FALSE"),                          // the TX and RX Reset FSMs must
           .RX_QPLL_USED             ("FALSE"),                          // share these two generic values
           .PHASE_ALIGNMENT_MANUAL   ("FALSE")                 // Decision if a manual phase-alignment is necessary or the automatic 
                                                                         // is enough. For single-lane applications the automatic alignment is 
                                                                         // sufficient              
             )     
gt7_rxresetfsm_i
             ( 
        .STABLE_CLOCK                   (SYSCLK_IN),
        .RXUSERCLK                      (GT7_RXUSRCLK_IN),
        .SOFT_RESET                     (SOFT_RESET_IN),
        .DONT_RESET_ON_DATA_ERROR       (DONT_RESET_ON_DATA_ERROR_IN),
        .QPLLREFCLKLOST                 (tied_to_ground_i),
        .CPLLREFCLKLOST                 (gt7_cpllrefclklost_i),
        .QPLLLOCK                       (tied_to_vcc_i),
        .CPLLLOCK                       (gt7_cplllock_i),
        .RXRESETDONE                    (gt7_rxresetdone_i),
        .MMCM_LOCK                      (tied_to_vcc_i),
        .RECCLK_STABLE                  (gt7_recclk_stable_i),
        .RECCLK_MONITOR_RESTART         (tied_to_ground_i),
        .DATA_VALID                     (GT7_DATA_VALID_IN),
        .TXUSERRDY                      (gt7_txuserrdy_i),
        .GTRXRESET                      (gt7_gtrxreset_t),
        .MMCM_RESET                     (),
        .QPLL_RESET                     (),
        .CPLL_RESET                     (),
        .RX_FSM_RESET_DONE              (GT7_RX_FSM_RESET_DONE_OUT),
        .RXUSERRDY                      (gt7_rxuserrdy_t),
        .RUN_PHALIGNMENT                (),
        .RESET_PHALIGNMENT              (),
        .PHALIGNMENT_DONE               (tied_to_vcc_i),
        .RXDFEAGCHOLD                   (gt7_rxdfeagchold_i),
        .RXDFELFHOLD                    (gt7_rxdfelfhold_i),
        .RXLPMLFHOLD                    (gt7_rxlpmlfhold_i),
        .RXLPMHFHOLD                    (gt7_rxlpmhfhold_i),
        .RETRY_COUNTER                  ()
           );

  always @(posedge SYSCLK_IN)
  begin
        if(gt0_gtrxreset_i)
        begin
          rx_cdrlocked       <= `DLY    1'b0;
          rx_cdrlock_counter <= `DLY    0;      
        end                
        else if (rx_cdrlock_counter == WAIT_TIME_CDRLOCK) 
        begin
          rx_cdrlocked       <= `DLY    1'b1;
          rx_cdrlock_counter <= `DLY    rx_cdrlock_counter;
        end
        else
          rx_cdrlock_counter <= `DLY    rx_cdrlock_counter + 1;
  end 

assign  gt0_recclk_stable_i                  =  rx_cdrlocked;
assign  gt1_recclk_stable_i                  =  rx_cdrlocked;
assign  gt2_recclk_stable_i                  =  rx_cdrlocked;
assign  gt3_recclk_stable_i                  =  rx_cdrlocked;
assign  gt4_recclk_stable_i                  =  rx_cdrlocked;
assign  gt5_recclk_stable_i                  =  rx_cdrlocked;
assign  gt6_recclk_stable_i                  =  rx_cdrlocked;
assign  gt7_recclk_stable_i                  =  rx_cdrlocked;








endmodule


